//Generate the verilog at 2024-10-31T21:13:53
module RVCPU (
clock,
io_interrupt,
io_master_arready,
io_master_arvalid,
io_master_awready,
io_master_awvalid,
io_master_bready,
io_master_bvalid,
io_master_rlast,
io_master_rready,
io_master_rvalid,
io_master_wlast,
io_master_wready,
io_master_wvalid,
io_slave_arready,
io_slave_arvalid,
io_slave_awready,
io_slave_awvalid,
io_slave_bready,
io_slave_bvalid,
io_slave_rlast,
io_slave_rready,
io_slave_rvalid,
io_slave_wlast,
io_slave_wready,
io_slave_wvalid,
reset,
io_master_araddr,
io_master_arburst,
io_master_arid,
io_master_arlen,
io_master_arsize,
io_master_awaddr,
io_master_awburst,
io_master_awid,
io_master_awlen,
io_master_awsize,
io_master_bid,
io_master_bresp,
io_master_rdata,
io_master_rid,
io_master_rresp,
io_master_wdata,
io_master_wstrb,
io_slave_araddr,
io_slave_arburst,
io_slave_arid,
io_slave_arlen,
io_slave_arsize,
io_slave_awaddr,
io_slave_awburst,
io_slave_awid,
io_slave_awlen,
io_slave_awsize,
io_slave_bid,
io_slave_bresp,
io_slave_rdata,
io_slave_rid,
io_slave_rresp,
io_slave_wdata,
io_slave_wstrb
);

input clock ;
input io_interrupt ;
input io_master_arready ;
output io_master_arvalid ;
input io_master_awready ;
output io_master_awvalid ;
output io_master_bready ;
input io_master_bvalid ;
input io_master_rlast ;
output io_master_rready ;
input io_master_rvalid ;
output io_master_wlast ;
input io_master_wready ;
output io_master_wvalid ;
output io_slave_arready ;
input io_slave_arvalid ;
output io_slave_awready ;
input io_slave_awvalid ;
input io_slave_bready ;
output io_slave_bvalid ;
output io_slave_rlast ;
input io_slave_rready ;
output io_slave_rvalid ;
input io_slave_wlast ;
output io_slave_wready ;
input io_slave_wvalid ;
input reset ;
output [31:0] io_master_araddr ;
output [1:0] io_master_arburst ;
output [3:0] io_master_arid ;
output [7:0] io_master_arlen ;
output [2:0] io_master_arsize ;
output [31:0] io_master_awaddr ;
output [1:0] io_master_awburst ;
output [3:0] io_master_awid ;
output [7:0] io_master_awlen ;
output [2:0] io_master_awsize ;
input [3:0] io_master_bid ;
input [1:0] io_master_bresp ;
input [31:0] io_master_rdata ;
input [3:0] io_master_rid ;
input [1:0] io_master_rresp ;
output [31:0] io_master_wdata ;
output [3:0] io_master_wstrb ;
input [31:0] io_slave_araddr ;
input [1:0] io_slave_arburst ;
input [3:0] io_slave_arid ;
input [7:0] io_slave_arlen ;
input [2:0] io_slave_arsize ;
input [31:0] io_slave_awaddr ;
input [1:0] io_slave_awburst ;
input [3:0] io_slave_awid ;
input [7:0] io_slave_awlen ;
input [2:0] io_slave_awsize ;
output [3:0] io_slave_bid ;
output [1:0] io_slave_bresp ;
output [31:0] io_slave_rdata ;
output [3:0] io_slave_rid ;
output [1:0] io_slave_rresp ;
input [31:0] io_slave_wdata ;
input [3:0] io_slave_wstrb ;

wire _00_ ;
wire _AXI4Interconnect_io_fanIn_0_arready ;
wire _AXI4Interconnect_io_fanIn_0_rvalid ;
wire _AXI4Interconnect_io_fanIn_1_arready ;
wire _AXI4Interconnect_io_fanIn_1_awready ;
wire _AXI4Interconnect_io_fanIn_1_bvalid ;
wire _AXI4Interconnect_io_fanIn_1_rvalid ;
wire _AXI4Interconnect_io_fanIn_1_wready ;
wire _AXI4Interconnect_io_fanOut_0_arvalid ;
wire _AXI4Interconnect_io_fanOut_0_awvalid ;
wire _AXI4Interconnect_io_fanOut_0_bready ;
wire _AXI4Interconnect_io_fanOut_0_rready ;
wire _AXI4Interconnect_io_fanOut_0_wvalid ;
wire _CLINT_io_arready ;
wire _CLINT_io_awready ;
wire _CLINT_io_bvalid ;
wire _CLINT_io_rvalid ;
wire _CLINT_io_wready ;
wire _EXU_io_LSUIn_bits_ren ;
wire _EXU_io_LSUIn_bits_wen ;
wire _EXU_io_LSUIn_valid ;
wire _EXU_io_LSUOut_ready ;
wire _EXU_io_in_ready ;
wire _EXU_io_out_bits_control_pcSrc ;
wire _EXU_io_out_bits_control_regWe ;
wire _EXU_io_out_valid ;
wire _IDU_io_in_ready ;
wire _IDU_io_out_bits_control_aluASrc ;
wire _IDU_io_out_bits_control_csrSrc ;
wire _IDU_io_out_bits_control_memRen ;
wire _IDU_io_out_bits_control_memWen ;
wire _IDU_io_out_bits_control_pcSrc ;
wire _IDU_io_out_bits_control_regWe ;
wire _IDU_io_out_valid ;
wire _IFU_io_in_ready ;
wire _IFU_io_master_arvalid ;
wire _IFU_io_master_rready ;
wire _IFU_io_out_valid ;
wire _LSU_io_in_ready ;
wire _LSU_io_master_arvalid ;
wire _LSU_io_master_awvalid ;
wire _LSU_io_master_bready ;
wire _LSU_io_master_rready ;
wire _LSU_io_master_wlast ;
wire _LSU_io_master_wvalid ;
wire _LSU_io_out_valid ;
wire _WBU_io_RegFileAccess_we ;
wire _WBU_io_in_ready ;
wire _WBU_io_out_valid ;
wire clock ;
wire io_interrupt ;
wire io_master_arready ;
wire io_master_arvalid ;
wire io_master_awready ;
wire io_master_awvalid ;
wire io_master_bready ;
wire io_master_bvalid ;
wire io_master_rlast ;
wire io_master_rready ;
wire io_master_rvalid ;
wire io_master_wlast ;
wire io_master_wready ;
wire io_master_wvalid ;
wire io_slave_arready ;
wire io_slave_arvalid ;
wire io_slave_awready ;
wire io_slave_awvalid ;
wire io_slave_bready ;
wire io_slave_bvalid ;
wire io_slave_rlast ;
wire io_slave_rready ;
wire io_slave_rvalid ;
wire io_slave_wlast ;
wire io_slave_wready ;
wire io_slave_wvalid ;
wire reset ;
wire \AXI4Interconnect/_0000_ ;
wire \AXI4Interconnect/_0001_ ;
wire \AXI4Interconnect/_0002_ ;
wire \AXI4Interconnect/_0003_ ;
wire \AXI4Interconnect/_0004_ ;
wire \AXI4Interconnect/_0005_ ;
wire \AXI4Interconnect/_0006_ ;
wire \AXI4Interconnect/_0007_ ;
wire \AXI4Interconnect/_0008_ ;
wire \AXI4Interconnect/_0009_ ;
wire \AXI4Interconnect/_0010_ ;
wire \AXI4Interconnect/_0011_ ;
wire \AXI4Interconnect/_0012_ ;
wire \AXI4Interconnect/_0013_ ;
wire \AXI4Interconnect/_0014_ ;
wire \AXI4Interconnect/_0015_ ;
wire \AXI4Interconnect/_0016_ ;
wire \AXI4Interconnect/_0017_ ;
wire \AXI4Interconnect/_0018_ ;
wire \AXI4Interconnect/_0019_ ;
wire \AXI4Interconnect/_0020_ ;
wire \AXI4Interconnect/_0021_ ;
wire \AXI4Interconnect/_0022_ ;
wire \AXI4Interconnect/_0023_ ;
wire \AXI4Interconnect/_0024_ ;
wire \AXI4Interconnect/_0025_ ;
wire \AXI4Interconnect/_0026_ ;
wire \AXI4Interconnect/_0027_ ;
wire \AXI4Interconnect/_0028_ ;
wire \AXI4Interconnect/_0029_ ;
wire \AXI4Interconnect/_0030_ ;
wire \AXI4Interconnect/_0031_ ;
wire \AXI4Interconnect/_0032_ ;
wire \AXI4Interconnect/_0033_ ;
wire \AXI4Interconnect/_0034_ ;
wire \AXI4Interconnect/_0035_ ;
wire \AXI4Interconnect/_0036_ ;
wire \AXI4Interconnect/_0037_ ;
wire \AXI4Interconnect/_0038_ ;
wire \AXI4Interconnect/_0039_ ;
wire \AXI4Interconnect/_0040_ ;
wire \AXI4Interconnect/_0041_ ;
wire \AXI4Interconnect/_0042_ ;
wire \AXI4Interconnect/_0043_ ;
wire \AXI4Interconnect/_0044_ ;
wire \AXI4Interconnect/_0045_ ;
wire \AXI4Interconnect/_0046_ ;
wire \AXI4Interconnect/_0047_ ;
wire \AXI4Interconnect/_0048_ ;
wire \AXI4Interconnect/_0049_ ;
wire \AXI4Interconnect/_0050_ ;
wire \AXI4Interconnect/_0051_ ;
wire \AXI4Interconnect/_0052_ ;
wire \AXI4Interconnect/_0053_ ;
wire \AXI4Interconnect/_0054_ ;
wire \AXI4Interconnect/_0055_ ;
wire \AXI4Interconnect/_0056_ ;
wire \AXI4Interconnect/_0057_ ;
wire \AXI4Interconnect/_0058_ ;
wire \AXI4Interconnect/_0059_ ;
wire \AXI4Interconnect/_0060_ ;
wire \AXI4Interconnect/_0061_ ;
wire \AXI4Interconnect/_0062_ ;
wire \AXI4Interconnect/_0063_ ;
wire \AXI4Interconnect/_0064_ ;
wire \AXI4Interconnect/_0065_ ;
wire \AXI4Interconnect/_0066_ ;
wire \AXI4Interconnect/_0067_ ;
wire \AXI4Interconnect/_0068_ ;
wire \AXI4Interconnect/_0069_ ;
wire \AXI4Interconnect/_0070_ ;
wire \AXI4Interconnect/_0071_ ;
wire \AXI4Interconnect/_0072_ ;
wire \AXI4Interconnect/_0073_ ;
wire \AXI4Interconnect/_0074_ ;
wire \AXI4Interconnect/_0075_ ;
wire \AXI4Interconnect/_0076_ ;
wire \AXI4Interconnect/_0077_ ;
wire \AXI4Interconnect/_0078_ ;
wire \AXI4Interconnect/_0079_ ;
wire \AXI4Interconnect/_0080_ ;
wire \AXI4Interconnect/_0081_ ;
wire \AXI4Interconnect/_0082_ ;
wire \AXI4Interconnect/_0083_ ;
wire \AXI4Interconnect/_0084_ ;
wire \AXI4Interconnect/_0085_ ;
wire \AXI4Interconnect/_0086_ ;
wire \AXI4Interconnect/_0087_ ;
wire \AXI4Interconnect/_0088_ ;
wire \AXI4Interconnect/_0089_ ;
wire \AXI4Interconnect/_0090_ ;
wire \AXI4Interconnect/_0091_ ;
wire \AXI4Interconnect/_0092_ ;
wire \AXI4Interconnect/_0093_ ;
wire \AXI4Interconnect/_0094_ ;
wire \AXI4Interconnect/_0095_ ;
wire \AXI4Interconnect/_0096_ ;
wire \AXI4Interconnect/_0097_ ;
wire \AXI4Interconnect/_0098_ ;
wire \AXI4Interconnect/_0099_ ;
wire \AXI4Interconnect/_0100_ ;
wire \AXI4Interconnect/_0101_ ;
wire \AXI4Interconnect/_0102_ ;
wire \AXI4Interconnect/_0103_ ;
wire \AXI4Interconnect/_0104_ ;
wire \AXI4Interconnect/_0105_ ;
wire \AXI4Interconnect/_0106_ ;
wire \AXI4Interconnect/_0107_ ;
wire \AXI4Interconnect/_0108_ ;
wire \AXI4Interconnect/_0109_ ;
wire \AXI4Interconnect/_0110_ ;
wire \AXI4Interconnect/_0111_ ;
wire \AXI4Interconnect/_0112_ ;
wire \AXI4Interconnect/_0113_ ;
wire \AXI4Interconnect/_0114_ ;
wire \AXI4Interconnect/_0115_ ;
wire \AXI4Interconnect/_0116_ ;
wire \AXI4Interconnect/_0117_ ;
wire \AXI4Interconnect/_0118_ ;
wire \AXI4Interconnect/_0119_ ;
wire \AXI4Interconnect/_0120_ ;
wire \AXI4Interconnect/_0121_ ;
wire \AXI4Interconnect/_0122_ ;
wire \AXI4Interconnect/_0123_ ;
wire \AXI4Interconnect/_0124_ ;
wire \AXI4Interconnect/_0125_ ;
wire \AXI4Interconnect/_0126_ ;
wire \AXI4Interconnect/_0127_ ;
wire \AXI4Interconnect/_0128_ ;
wire \AXI4Interconnect/_0129_ ;
wire \AXI4Interconnect/_0130_ ;
wire \AXI4Interconnect/_0131_ ;
wire \AXI4Interconnect/_0132_ ;
wire \AXI4Interconnect/_0133_ ;
wire \AXI4Interconnect/_0134_ ;
wire \AXI4Interconnect/_0135_ ;
wire \AXI4Interconnect/_0136_ ;
wire \AXI4Interconnect/_0137_ ;
wire \AXI4Interconnect/_0138_ ;
wire \AXI4Interconnect/_0139_ ;
wire \AXI4Interconnect/_0140_ ;
wire \AXI4Interconnect/_0141_ ;
wire \AXI4Interconnect/_0142_ ;
wire \AXI4Interconnect/_0143_ ;
wire \AXI4Interconnect/_0144_ ;
wire \AXI4Interconnect/_0145_ ;
wire \AXI4Interconnect/_0146_ ;
wire \AXI4Interconnect/_0147_ ;
wire \AXI4Interconnect/_0148_ ;
wire \AXI4Interconnect/_0149_ ;
wire \AXI4Interconnect/_0150_ ;
wire \AXI4Interconnect/_0151_ ;
wire \AXI4Interconnect/_0152_ ;
wire \AXI4Interconnect/_0153_ ;
wire \AXI4Interconnect/_0154_ ;
wire \AXI4Interconnect/_0155_ ;
wire \AXI4Interconnect/_0156_ ;
wire \AXI4Interconnect/_0157_ ;
wire \AXI4Interconnect/_0158_ ;
wire \AXI4Interconnect/_0159_ ;
wire \AXI4Interconnect/_0160_ ;
wire \AXI4Interconnect/_0161_ ;
wire \AXI4Interconnect/_0162_ ;
wire \AXI4Interconnect/_0163_ ;
wire \AXI4Interconnect/_0164_ ;
wire \AXI4Interconnect/_0165_ ;
wire \AXI4Interconnect/_0166_ ;
wire \AXI4Interconnect/_0167_ ;
wire \AXI4Interconnect/_0168_ ;
wire \AXI4Interconnect/_0169_ ;
wire \AXI4Interconnect/_0170_ ;
wire \AXI4Interconnect/_0171_ ;
wire \AXI4Interconnect/_0172_ ;
wire \AXI4Interconnect/_0173_ ;
wire \AXI4Interconnect/_0174_ ;
wire \AXI4Interconnect/_0175_ ;
wire \AXI4Interconnect/_0176_ ;
wire \AXI4Interconnect/_0177_ ;
wire \AXI4Interconnect/_0178_ ;
wire \AXI4Interconnect/_0179_ ;
wire \AXI4Interconnect/_0180_ ;
wire \AXI4Interconnect/_0181_ ;
wire \AXI4Interconnect/_0182_ ;
wire \AXI4Interconnect/_0183_ ;
wire \AXI4Interconnect/_0184_ ;
wire \AXI4Interconnect/_0185_ ;
wire \AXI4Interconnect/_0186_ ;
wire \AXI4Interconnect/_0187_ ;
wire \AXI4Interconnect/_0188_ ;
wire \AXI4Interconnect/_0189_ ;
wire \AXI4Interconnect/_0190_ ;
wire \AXI4Interconnect/_0191_ ;
wire \AXI4Interconnect/_0192_ ;
wire \AXI4Interconnect/_0193_ ;
wire \AXI4Interconnect/_0194_ ;
wire \AXI4Interconnect/_0195_ ;
wire \AXI4Interconnect/_0196_ ;
wire \AXI4Interconnect/_0197_ ;
wire \AXI4Interconnect/_0198_ ;
wire \AXI4Interconnect/_0199_ ;
wire \AXI4Interconnect/_0200_ ;
wire \AXI4Interconnect/_0201_ ;
wire \AXI4Interconnect/_0202_ ;
wire \AXI4Interconnect/_0203_ ;
wire \AXI4Interconnect/_0204_ ;
wire \AXI4Interconnect/_0205_ ;
wire \AXI4Interconnect/_0206_ ;
wire \AXI4Interconnect/_0207_ ;
wire \AXI4Interconnect/_0208_ ;
wire \AXI4Interconnect/_0209_ ;
wire \AXI4Interconnect/_0210_ ;
wire \AXI4Interconnect/_0211_ ;
wire \AXI4Interconnect/_0212_ ;
wire \AXI4Interconnect/_0213_ ;
wire \AXI4Interconnect/_0214_ ;
wire \AXI4Interconnect/_0215_ ;
wire \AXI4Interconnect/_0216_ ;
wire \AXI4Interconnect/_0217_ ;
wire \AXI4Interconnect/_0218_ ;
wire \AXI4Interconnect/_0219_ ;
wire \AXI4Interconnect/_0220_ ;
wire \AXI4Interconnect/_0221_ ;
wire \AXI4Interconnect/_0222_ ;
wire \AXI4Interconnect/_0223_ ;
wire \AXI4Interconnect/_0224_ ;
wire \AXI4Interconnect/_0225_ ;
wire \AXI4Interconnect/_0226_ ;
wire \AXI4Interconnect/_0227_ ;
wire \AXI4Interconnect/_0228_ ;
wire \AXI4Interconnect/_0229_ ;
wire \AXI4Interconnect/_0230_ ;
wire \AXI4Interconnect/_0231_ ;
wire \AXI4Interconnect/_0232_ ;
wire \AXI4Interconnect/_0233_ ;
wire \AXI4Interconnect/_0234_ ;
wire \AXI4Interconnect/_0235_ ;
wire \AXI4Interconnect/_0236_ ;
wire \AXI4Interconnect/_0237_ ;
wire \AXI4Interconnect/_0238_ ;
wire \AXI4Interconnect/_0239_ ;
wire \AXI4Interconnect/_0240_ ;
wire \AXI4Interconnect/_0241_ ;
wire \AXI4Interconnect/_0242_ ;
wire \AXI4Interconnect/_0243_ ;
wire \AXI4Interconnect/_0244_ ;
wire \AXI4Interconnect/_0245_ ;
wire \AXI4Interconnect/_0246_ ;
wire \AXI4Interconnect/_0247_ ;
wire \AXI4Interconnect/_0248_ ;
wire \AXI4Interconnect/_0249_ ;
wire \AXI4Interconnect/_0250_ ;
wire \AXI4Interconnect/_0251_ ;
wire \AXI4Interconnect/_0252_ ;
wire \AXI4Interconnect/_0253_ ;
wire \AXI4Interconnect/_0254_ ;
wire \AXI4Interconnect/_0255_ ;
wire \AXI4Interconnect/_0256_ ;
wire \AXI4Interconnect/_0257_ ;
wire \AXI4Interconnect/_0258_ ;
wire \AXI4Interconnect/_0259_ ;
wire \AXI4Interconnect/_0260_ ;
wire \AXI4Interconnect/_0261_ ;
wire \AXI4Interconnect/_0262_ ;
wire \AXI4Interconnect/_0263_ ;
wire \AXI4Interconnect/_0264_ ;
wire \AXI4Interconnect/_0265_ ;
wire \AXI4Interconnect/_0266_ ;
wire \AXI4Interconnect/_0267_ ;
wire \AXI4Interconnect/_0268_ ;
wire \AXI4Interconnect/_0269_ ;
wire \AXI4Interconnect/_0270_ ;
wire \AXI4Interconnect/_0271_ ;
wire \AXI4Interconnect/_0272_ ;
wire \AXI4Interconnect/_0273_ ;
wire \AXI4Interconnect/_0274_ ;
wire \AXI4Interconnect/_0275_ ;
wire \AXI4Interconnect/_0276_ ;
wire \AXI4Interconnect/_0277_ ;
wire \AXI4Interconnect/_0278_ ;
wire \AXI4Interconnect/_0279_ ;
wire \AXI4Interconnect/_0280_ ;
wire \AXI4Interconnect/_0281_ ;
wire \AXI4Interconnect/_0282_ ;
wire \AXI4Interconnect/_0283_ ;
wire \AXI4Interconnect/_0284_ ;
wire \AXI4Interconnect/_0285_ ;
wire \AXI4Interconnect/_0286_ ;
wire \AXI4Interconnect/_0287_ ;
wire \AXI4Interconnect/_0288_ ;
wire \AXI4Interconnect/_0289_ ;
wire \AXI4Interconnect/_0290_ ;
wire \AXI4Interconnect/_0291_ ;
wire \AXI4Interconnect/_0292_ ;
wire \AXI4Interconnect/_0293_ ;
wire \AXI4Interconnect/_0294_ ;
wire \AXI4Interconnect/_0295_ ;
wire \AXI4Interconnect/_0296_ ;
wire \AXI4Interconnect/_0297_ ;
wire \AXI4Interconnect/_0298_ ;
wire \AXI4Interconnect/_0299_ ;
wire \AXI4Interconnect/_0300_ ;
wire \AXI4Interconnect/_0301_ ;
wire \AXI4Interconnect/_0302_ ;
wire \AXI4Interconnect/_0303_ ;
wire \AXI4Interconnect/_0304_ ;
wire \AXI4Interconnect/_0305_ ;
wire \AXI4Interconnect/_0306_ ;
wire \AXI4Interconnect/_0307_ ;
wire \AXI4Interconnect/_0308_ ;
wire \AXI4Interconnect/_0309_ ;
wire \AXI4Interconnect/_0310_ ;
wire \AXI4Interconnect/_0311_ ;
wire \AXI4Interconnect/_0312_ ;
wire \AXI4Interconnect/_0313_ ;
wire \AXI4Interconnect/_0314_ ;
wire \AXI4Interconnect/_0315_ ;
wire \AXI4Interconnect/_0316_ ;
wire \AXI4Interconnect/_0317_ ;
wire \AXI4Interconnect/_0318_ ;
wire \AXI4Interconnect/_0319_ ;
wire \AXI4Interconnect/_0320_ ;
wire \AXI4Interconnect/_0321_ ;
wire \AXI4Interconnect/_0322_ ;
wire \AXI4Interconnect/_0323_ ;
wire \AXI4Interconnect/_0324_ ;
wire \AXI4Interconnect/_0325_ ;
wire \AXI4Interconnect/_0326_ ;
wire \AXI4Interconnect/_0327_ ;
wire \AXI4Interconnect/_0328_ ;
wire \AXI4Interconnect/_0329_ ;
wire \AXI4Interconnect/_0330_ ;
wire \AXI4Interconnect/_0331_ ;
wire \AXI4Interconnect/_0332_ ;
wire \AXI4Interconnect/_0333_ ;
wire \AXI4Interconnect/_0334_ ;
wire \AXI4Interconnect/_0335_ ;
wire \AXI4Interconnect/_0336_ ;
wire \AXI4Interconnect/_0337_ ;
wire \AXI4Interconnect/_0338_ ;
wire \AXI4Interconnect/_0339_ ;
wire \AXI4Interconnect/_0340_ ;
wire \AXI4Interconnect/_0341_ ;
wire \AXI4Interconnect/_0342_ ;
wire \AXI4Interconnect/_0343_ ;
wire \AXI4Interconnect/_0344_ ;
wire \AXI4Interconnect/_0345_ ;
wire \AXI4Interconnect/_0346_ ;
wire \AXI4Interconnect/_0347_ ;
wire \AXI4Interconnect/_0348_ ;
wire \AXI4Interconnect/_0349_ ;
wire \AXI4Interconnect/_0350_ ;
wire \AXI4Interconnect/_0351_ ;
wire \AXI4Interconnect/_0352_ ;
wire \AXI4Interconnect/_0353_ ;
wire \AXI4Interconnect/_0354_ ;
wire \AXI4Interconnect/_0355_ ;
wire \AXI4Interconnect/_0356_ ;
wire \AXI4Interconnect/_0357_ ;
wire \AXI4Interconnect/_0358_ ;
wire \AXI4Interconnect/_0359_ ;
wire \AXI4Interconnect/_0360_ ;
wire \AXI4Interconnect/_0361_ ;
wire \AXI4Interconnect/_0362_ ;
wire \AXI4Interconnect/_0363_ ;
wire \AXI4Interconnect/_0364_ ;
wire \AXI4Interconnect/_0365_ ;
wire \AXI4Interconnect/_0366_ ;
wire \AXI4Interconnect/_0367_ ;
wire \AXI4Interconnect/_0368_ ;
wire \AXI4Interconnect/_0369_ ;
wire \AXI4Interconnect/_0370_ ;
wire \AXI4Interconnect/_0371_ ;
wire \AXI4Interconnect/_0372_ ;
wire \AXI4Interconnect/_0373_ ;
wire \AXI4Interconnect/_0374_ ;
wire \AXI4Interconnect/_0375_ ;
wire \AXI4Interconnect/_0376_ ;
wire \AXI4Interconnect/_0377_ ;
wire \AXI4Interconnect/_0378_ ;
wire \AXI4Interconnect/_0379_ ;
wire \AXI4Interconnect/_0380_ ;
wire \AXI4Interconnect/_0381_ ;
wire \AXI4Interconnect/_0382_ ;
wire \AXI4Interconnect/_0383_ ;
wire \AXI4Interconnect/_0384_ ;
wire \AXI4Interconnect/_0385_ ;
wire \AXI4Interconnect/_0386_ ;
wire \AXI4Interconnect/_0387_ ;
wire \AXI4Interconnect/_0388_ ;
wire \AXI4Interconnect/_0389_ ;
wire \AXI4Interconnect/_0390_ ;
wire \AXI4Interconnect/_0391_ ;
wire \AXI4Interconnect/_0392_ ;
wire \AXI4Interconnect/_0393_ ;
wire \AXI4Interconnect/_0394_ ;
wire \AXI4Interconnect/_0395_ ;
wire \AXI4Interconnect/_0396_ ;
wire \AXI4Interconnect/_0397_ ;
wire \AXI4Interconnect/_0398_ ;
wire \AXI4Interconnect/_0399_ ;
wire \AXI4Interconnect/_0400_ ;
wire \AXI4Interconnect/_0401_ ;
wire \AXI4Interconnect/_0402_ ;
wire \AXI4Interconnect/_0403_ ;
wire \AXI4Interconnect/_0404_ ;
wire \AXI4Interconnect/_0405_ ;
wire \AXI4Interconnect/_0406_ ;
wire \AXI4Interconnect/_0407_ ;
wire \AXI4Interconnect/_0408_ ;
wire \AXI4Interconnect/_0409_ ;
wire \AXI4Interconnect/_0410_ ;
wire \AXI4Interconnect/_0411_ ;
wire \AXI4Interconnect/_0412_ ;
wire \AXI4Interconnect/_0413_ ;
wire \AXI4Interconnect/_0414_ ;
wire \AXI4Interconnect/_0415_ ;
wire \AXI4Interconnect/_0416_ ;
wire \AXI4Interconnect/_0417_ ;
wire \AXI4Interconnect/_0418_ ;
wire \AXI4Interconnect/_0419_ ;
wire \AXI4Interconnect/_0420_ ;
wire \AXI4Interconnect/_0421_ ;
wire \AXI4Interconnect/_0422_ ;
wire \AXI4Interconnect/_0423_ ;
wire \AXI4Interconnect/_0424_ ;
wire \AXI4Interconnect/_0425_ ;
wire \AXI4Interconnect/_0426_ ;
wire \AXI4Interconnect/_0427_ ;
wire \AXI4Interconnect/_0428_ ;
wire \AXI4Interconnect/_0429_ ;
wire \AXI4Interconnect/_0430_ ;
wire \AXI4Interconnect/_0431_ ;
wire \AXI4Interconnect/_0432_ ;
wire \AXI4Interconnect/_0433_ ;
wire \AXI4Interconnect/_0434_ ;
wire \AXI4Interconnect/_0435_ ;
wire \AXI4Interconnect/_0436_ ;
wire \AXI4Interconnect/_0437_ ;
wire \AXI4Interconnect/_0438_ ;
wire \AXI4Interconnect/_0439_ ;
wire \AXI4Interconnect/_0440_ ;
wire \AXI4Interconnect/_0441_ ;
wire \AXI4Interconnect/_0442_ ;
wire \AXI4Interconnect/_0443_ ;
wire \AXI4Interconnect/_0444_ ;
wire \AXI4Interconnect/_0445_ ;
wire \AXI4Interconnect/_0446_ ;
wire \AXI4Interconnect/_0447_ ;
wire \AXI4Interconnect/_0448_ ;
wire \AXI4Interconnect/_0449_ ;
wire \AXI4Interconnect/_0450_ ;
wire \AXI4Interconnect/_0451_ ;
wire \AXI4Interconnect/_0452_ ;
wire \AXI4Interconnect/_0453_ ;
wire \AXI4Interconnect/_0454_ ;
wire \AXI4Interconnect/_0455_ ;
wire \AXI4Interconnect/_0456_ ;
wire \AXI4Interconnect/_0457_ ;
wire \AXI4Interconnect/_0458_ ;
wire \AXI4Interconnect/_0459_ ;
wire \AXI4Interconnect/_0460_ ;
wire \AXI4Interconnect/_0461_ ;
wire \AXI4Interconnect/_0462_ ;
wire \AXI4Interconnect/_0463_ ;
wire \AXI4Interconnect/_0464_ ;
wire \AXI4Interconnect/_0465_ ;
wire \AXI4Interconnect/_0466_ ;
wire \AXI4Interconnect/_0467_ ;
wire \AXI4Interconnect/_0468_ ;
wire \AXI4Interconnect/_0469_ ;
wire \AXI4Interconnect/_0470_ ;
wire \AXI4Interconnect/_0471_ ;
wire \AXI4Interconnect/_0472_ ;
wire \AXI4Interconnect/_0473_ ;
wire \AXI4Interconnect/_0474_ ;
wire \AXI4Interconnect/_0475_ ;
wire \AXI4Interconnect/_0476_ ;
wire \AXI4Interconnect/_0477_ ;
wire \AXI4Interconnect/_0478_ ;
wire \AXI4Interconnect/_0479_ ;
wire \AXI4Interconnect/_0480_ ;
wire \AXI4Interconnect/_0481_ ;
wire \AXI4Interconnect/_0482_ ;
wire \AXI4Interconnect/_0483_ ;
wire \AXI4Interconnect/_0484_ ;
wire \AXI4Interconnect/_0485_ ;
wire \AXI4Interconnect/_0486_ ;
wire \AXI4Interconnect/_0487_ ;
wire \AXI4Interconnect/_0488_ ;
wire \AXI4Interconnect/_0489_ ;
wire \AXI4Interconnect/_0490_ ;
wire \AXI4Interconnect/_0491_ ;
wire \AXI4Interconnect/_0492_ ;
wire \AXI4Interconnect/_0493_ ;
wire \AXI4Interconnect/_0494_ ;
wire \AXI4Interconnect/_0495_ ;
wire \AXI4Interconnect/_0496_ ;
wire \AXI4Interconnect/_0497_ ;
wire \AXI4Interconnect/_0498_ ;
wire \AXI4Interconnect/_0499_ ;
wire \AXI4Interconnect/_0500_ ;
wire \AXI4Interconnect/_0501_ ;
wire \AXI4Interconnect/_0502_ ;
wire \AXI4Interconnect/_0503_ ;
wire \AXI4Interconnect/_0504_ ;
wire \AXI4Interconnect/_0505_ ;
wire \AXI4Interconnect/_0506_ ;
wire \AXI4Interconnect/_0507_ ;
wire \AXI4Interconnect/_0508_ ;
wire \AXI4Interconnect/_0509_ ;
wire \AXI4Interconnect/_0510_ ;
wire \AXI4Interconnect/_0511_ ;
wire \AXI4Interconnect/_0512_ ;
wire \AXI4Interconnect/_0513_ ;
wire \AXI4Interconnect/_0514_ ;
wire \AXI4Interconnect/_0515_ ;
wire \AXI4Interconnect/_0516_ ;
wire \AXI4Interconnect/_0517_ ;
wire \AXI4Interconnect/_0518_ ;
wire \AXI4Interconnect/_0519_ ;
wire \AXI4Interconnect/_0520_ ;
wire \AXI4Interconnect/_0521_ ;
wire \AXI4Interconnect/_0522_ ;
wire \AXI4Interconnect/_0523_ ;
wire \AXI4Interconnect/_0524_ ;
wire \AXI4Interconnect/_0525_ ;
wire \AXI4Interconnect/_0526_ ;
wire \AXI4Interconnect/_0527_ ;
wire \AXI4Interconnect/_0528_ ;
wire \AXI4Interconnect/_0529_ ;
wire \AXI4Interconnect/_0530_ ;
wire \AXI4Interconnect/_0531_ ;
wire \AXI4Interconnect/_0532_ ;
wire \AXI4Interconnect/_0533_ ;
wire \AXI4Interconnect/_0534_ ;
wire \AXI4Interconnect/_0535_ ;
wire \AXI4Interconnect/_0536_ ;
wire \AXI4Interconnect/_0537_ ;
wire \AXI4Interconnect/_0538_ ;
wire \AXI4Interconnect/_0539_ ;
wire \AXI4Interconnect/_0540_ ;
wire \AXI4Interconnect/_0541_ ;
wire \AXI4Interconnect/_0542_ ;
wire \AXI4Interconnect/_0543_ ;
wire \AXI4Interconnect/_0544_ ;
wire \AXI4Interconnect/_0545_ ;
wire \AXI4Interconnect/_0546_ ;
wire \AXI4Interconnect/_0547_ ;
wire \AXI4Interconnect/_0548_ ;
wire \AXI4Interconnect/_0549_ ;
wire \AXI4Interconnect/_0550_ ;
wire \AXI4Interconnect/_0551_ ;
wire \AXI4Interconnect/_0552_ ;
wire \AXI4Interconnect/_0553_ ;
wire \AXI4Interconnect/_0554_ ;
wire \AXI4Interconnect/_0555_ ;
wire \AXI4Interconnect/_0556_ ;
wire \AXI4Interconnect/_0557_ ;
wire \AXI4Interconnect/_0558_ ;
wire \AXI4Interconnect/_0559_ ;
wire \AXI4Interconnect/_0560_ ;
wire \AXI4Interconnect/_0561_ ;
wire \AXI4Interconnect/_0562_ ;
wire \AXI4Interconnect/_0563_ ;
wire \AXI4Interconnect/_0564_ ;
wire \AXI4Interconnect/_0565_ ;
wire \AXI4Interconnect/_0566_ ;
wire \AXI4Interconnect/_0567_ ;
wire \AXI4Interconnect/_0568_ ;
wire \AXI4Interconnect/_0569_ ;
wire \AXI4Interconnect/_0570_ ;
wire \AXI4Interconnect/_0571_ ;
wire \AXI4Interconnect/_0572_ ;
wire \AXI4Interconnect/_0573_ ;
wire \AXI4Interconnect/_0574_ ;
wire \AXI4Interconnect/_0575_ ;
wire \AXI4Interconnect/_0576_ ;
wire \AXI4Interconnect/_0577_ ;
wire \AXI4Interconnect/_0578_ ;
wire \AXI4Interconnect/_0579_ ;
wire \AXI4Interconnect/_0580_ ;
wire \AXI4Interconnect/_0581_ ;
wire \AXI4Interconnect/_0582_ ;
wire \AXI4Interconnect/_0583_ ;
wire \AXI4Interconnect/_0584_ ;
wire \AXI4Interconnect/_0585_ ;
wire \AXI4Interconnect/_0586_ ;
wire \AXI4Interconnect/_0587_ ;
wire \AXI4Interconnect/_0588_ ;
wire \AXI4Interconnect/_0589_ ;
wire \AXI4Interconnect/_0590_ ;
wire \AXI4Interconnect/_0591_ ;
wire \AXI4Interconnect/_0592_ ;
wire \AXI4Interconnect/_0593_ ;
wire \AXI4Interconnect/_0594_ ;
wire \AXI4Interconnect/_0595_ ;
wire \AXI4Interconnect/_0596_ ;
wire \AXI4Interconnect/_0597_ ;
wire \AXI4Interconnect/_0598_ ;
wire \AXI4Interconnect/_0599_ ;
wire \AXI4Interconnect/_0600_ ;
wire \AXI4Interconnect/_0601_ ;
wire \AXI4Interconnect/_0602_ ;
wire \AXI4Interconnect/_0603_ ;
wire \AXI4Interconnect/_0604_ ;
wire \AXI4Interconnect/_0605_ ;
wire \AXI4Interconnect/_0606_ ;
wire \AXI4Interconnect/_0607_ ;
wire \AXI4Interconnect/_0608_ ;
wire \AXI4Interconnect/_0609_ ;
wire \AXI4Interconnect/_0610_ ;
wire \AXI4Interconnect/_0611_ ;
wire \AXI4Interconnect/_0612_ ;
wire \AXI4Interconnect/_0613_ ;
wire \AXI4Interconnect/_0614_ ;
wire \AXI4Interconnect/_0615_ ;
wire \AXI4Interconnect/_0616_ ;
wire \AXI4Interconnect/_0617_ ;
wire \AXI4Interconnect/_0618_ ;
wire \AXI4Interconnect/_0619_ ;
wire \AXI4Interconnect/_0620_ ;
wire \AXI4Interconnect/_0621_ ;
wire \AXI4Interconnect/_0622_ ;
wire \AXI4Interconnect/_0623_ ;
wire \AXI4Interconnect/_0624_ ;
wire \AXI4Interconnect/_0625_ ;
wire \AXI4Interconnect/_0626_ ;
wire \AXI4Interconnect/_0627_ ;
wire \AXI4Interconnect/_0628_ ;
wire \AXI4Interconnect/_0629_ ;
wire \AXI4Interconnect/_0630_ ;
wire \AXI4Interconnect/_0631_ ;
wire \AXI4Interconnect/_0632_ ;
wire \AXI4Interconnect/_0633_ ;
wire \AXI4Interconnect/_0634_ ;
wire \AXI4Interconnect/_0635_ ;
wire \AXI4Interconnect/_0636_ ;
wire \AXI4Interconnect/_0637_ ;
wire \AXI4Interconnect/_0638_ ;
wire \AXI4Interconnect/_0639_ ;
wire \AXI4Interconnect/_0640_ ;
wire \AXI4Interconnect/_0641_ ;
wire \AXI4Interconnect/_0642_ ;
wire \AXI4Interconnect/_0643_ ;
wire \AXI4Interconnect/_0644_ ;
wire \AXI4Interconnect/_0645_ ;
wire \AXI4Interconnect/_0646_ ;
wire \AXI4Interconnect/_0647_ ;
wire \AXI4Interconnect/_0648_ ;
wire \AXI4Interconnect/_0649_ ;
wire \AXI4Interconnect/_0650_ ;
wire \AXI4Interconnect/_0651_ ;
wire \AXI4Interconnect/_0652_ ;
wire \AXI4Interconnect/_0653_ ;
wire \AXI4Interconnect/_0654_ ;
wire \AXI4Interconnect/_0655_ ;
wire \AXI4Interconnect/_0656_ ;
wire \AXI4Interconnect/_0657_ ;
wire \AXI4Interconnect/_0658_ ;
wire \AXI4Interconnect/_0659_ ;
wire \AXI4Interconnect/_0660_ ;
wire \AXI4Interconnect/_0661_ ;
wire \AXI4Interconnect/_0662_ ;
wire \AXI4Interconnect/_0663_ ;
wire \AXI4Interconnect/_0664_ ;
wire \AXI4Interconnect/_0665_ ;
wire \AXI4Interconnect/_0666_ ;
wire \AXI4Interconnect/_0667_ ;
wire \AXI4Interconnect/_0668_ ;
wire \AXI4Interconnect/_0669_ ;
wire \AXI4Interconnect/_0670_ ;
wire \AXI4Interconnect/_0671_ ;
wire \AXI4Interconnect/_0672_ ;
wire \AXI4Interconnect/_0673_ ;
wire \AXI4Interconnect/_0674_ ;
wire \AXI4Interconnect/_0675_ ;
wire \AXI4Interconnect/_0676_ ;
wire \AXI4Interconnect/_0677_ ;
wire \AXI4Interconnect/_0678_ ;
wire \AXI4Interconnect/_0679_ ;
wire \AXI4Interconnect/_0680_ ;
wire \AXI4Interconnect/_0681_ ;
wire \AXI4Interconnect/_0682_ ;
wire \AXI4Interconnect/_0683_ ;
wire \AXI4Interconnect/_0684_ ;
wire \AXI4Interconnect/_0685_ ;
wire \AXI4Interconnect/_0686_ ;
wire \AXI4Interconnect/_0687_ ;
wire \AXI4Interconnect/_0688_ ;
wire \AXI4Interconnect/_0689_ ;
wire \AXI4Interconnect/_0690_ ;
wire \AXI4Interconnect/_0691_ ;
wire \AXI4Interconnect/_0692_ ;
wire \AXI4Interconnect/_0693_ ;
wire \AXI4Interconnect/_0694_ ;
wire \AXI4Interconnect/_0695_ ;
wire \AXI4Interconnect/_0696_ ;
wire \AXI4Interconnect/_0697_ ;
wire \AXI4Interconnect/_0698_ ;
wire \AXI4Interconnect/_0699_ ;
wire \AXI4Interconnect/_0700_ ;
wire \AXI4Interconnect/_0701_ ;
wire \AXI4Interconnect/_0702_ ;
wire \AXI4Interconnect/_0703_ ;
wire \AXI4Interconnect/_0704_ ;
wire \AXI4Interconnect/_0705_ ;
wire \AXI4Interconnect/_0706_ ;
wire \AXI4Interconnect/_0707_ ;
wire \AXI4Interconnect/_0708_ ;
wire \AXI4Interconnect/_0709_ ;
wire \AXI4Interconnect/_0710_ ;
wire \AXI4Interconnect/_0711_ ;
wire \AXI4Interconnect/_0712_ ;
wire \AXI4Interconnect/_0713_ ;
wire \AXI4Interconnect/_0714_ ;
wire \AXI4Interconnect/_0715_ ;
wire \AXI4Interconnect/_0716_ ;
wire \AXI4Interconnect/_0717_ ;
wire \AXI4Interconnect/_0718_ ;
wire \AXI4Interconnect/_0719_ ;
wire \AXI4Interconnect/_0720_ ;
wire \AXI4Interconnect/_0721_ ;
wire \AXI4Interconnect/_0722_ ;
wire \AXI4Interconnect/_0723_ ;
wire \AXI4Interconnect/_0724_ ;
wire \AXI4Interconnect/_0725_ ;
wire \AXI4Interconnect/_0726_ ;
wire \AXI4Interconnect/_0727_ ;
wire \AXI4Interconnect/_0728_ ;
wire \AXI4Interconnect/_0729_ ;
wire \AXI4Interconnect/_0730_ ;
wire \AXI4Interconnect/_0731_ ;
wire \AXI4Interconnect/_0732_ ;
wire \AXI4Interconnect/_0733_ ;
wire \AXI4Interconnect/_0734_ ;
wire \AXI4Interconnect/_0735_ ;
wire \AXI4Interconnect/_0736_ ;
wire \AXI4Interconnect/_0737_ ;
wire \AXI4Interconnect/_0738_ ;
wire \AXI4Interconnect/_0739_ ;
wire \AXI4Interconnect/_0740_ ;
wire \AXI4Interconnect/_0741_ ;
wire \AXI4Interconnect/_0742_ ;
wire \AXI4Interconnect/_0743_ ;
wire \AXI4Interconnect/_0744_ ;
wire \AXI4Interconnect/_0745_ ;
wire \AXI4Interconnect/_0746_ ;
wire \AXI4Interconnect/_0747_ ;
wire \AXI4Interconnect/_0748_ ;
wire \AXI4Interconnect/_0749_ ;
wire \AXI4Interconnect/_0750_ ;
wire \AXI4Interconnect/_0751_ ;
wire \AXI4Interconnect/_0752_ ;
wire \AXI4Interconnect/_0753_ ;
wire \AXI4Interconnect/_0754_ ;
wire \AXI4Interconnect/_0755_ ;
wire \AXI4Interconnect/_0756_ ;
wire \AXI4Interconnect/_0757_ ;
wire \AXI4Interconnect/_0758_ ;
wire \AXI4Interconnect/_0759_ ;
wire \AXI4Interconnect/_0760_ ;
wire \AXI4Interconnect/_0761_ ;
wire \AXI4Interconnect/_0762_ ;
wire \AXI4Interconnect/_0763_ ;
wire \AXI4Interconnect/_0764_ ;
wire \AXI4Interconnect/_0765_ ;
wire \AXI4Interconnect/_0766_ ;
wire \AXI4Interconnect/_0767_ ;
wire \AXI4Interconnect/_0768_ ;
wire \AXI4Interconnect/_0769_ ;
wire \AXI4Interconnect/_0770_ ;
wire \AXI4Interconnect/_0771_ ;
wire \AXI4Interconnect/_0772_ ;
wire \AXI4Interconnect/_0773_ ;
wire \AXI4Interconnect/_0774_ ;
wire \AXI4Interconnect/_0775_ ;
wire \AXI4Interconnect/_0776_ ;
wire \AXI4Interconnect/_0777_ ;
wire \AXI4Interconnect/_0778_ ;
wire \AXI4Interconnect/_0779_ ;
wire \AXI4Interconnect/_0780_ ;
wire \AXI4Interconnect/_0781_ ;
wire \AXI4Interconnect/_0782_ ;
wire \AXI4Interconnect/_0783_ ;
wire \AXI4Interconnect/_0784_ ;
wire \AXI4Interconnect/_0785_ ;
wire \AXI4Interconnect/_0786_ ;
wire \AXI4Interconnect/_0787_ ;
wire \AXI4Interconnect/_0788_ ;
wire \AXI4Interconnect/_0789_ ;
wire \AXI4Interconnect/_0790_ ;
wire \AXI4Interconnect/_0791_ ;
wire \AXI4Interconnect/_0792_ ;
wire \AXI4Interconnect/_0793_ ;
wire \AXI4Interconnect/_0794_ ;
wire \AXI4Interconnect/_0795_ ;
wire \AXI4Interconnect/_0796_ ;
wire \AXI4Interconnect/_0797_ ;
wire \AXI4Interconnect/_0798_ ;
wire \AXI4Interconnect/_0799_ ;
wire \AXI4Interconnect/_0800_ ;
wire \AXI4Interconnect/_0801_ ;
wire \AXI4Interconnect/_0802_ ;
wire \AXI4Interconnect/_0803_ ;
wire \AXI4Interconnect/_0804_ ;
wire \AXI4Interconnect/_0805_ ;
wire \AXI4Interconnect/_0806_ ;
wire \AXI4Interconnect/_0807_ ;
wire \AXI4Interconnect/_0808_ ;
wire \AXI4Interconnect/_0809_ ;
wire \AXI4Interconnect/_0810_ ;
wire \AXI4Interconnect/_0811_ ;
wire \AXI4Interconnect/_0812_ ;
wire \AXI4Interconnect/_0813_ ;
wire \AXI4Interconnect/_0814_ ;
wire \AXI4Interconnect/_0815_ ;
wire \AXI4Interconnect/_0816_ ;
wire \AXI4Interconnect/_0817_ ;
wire \AXI4Interconnect/_0818_ ;
wire \AXI4Interconnect/_0819_ ;
wire \AXI4Interconnect/_0820_ ;
wire \AXI4Interconnect/_0821_ ;
wire \AXI4Interconnect/_0822_ ;
wire \AXI4Interconnect/_0823_ ;
wire \AXI4Interconnect/_0824_ ;
wire \AXI4Interconnect/_0825_ ;
wire \AXI4Interconnect/_0826_ ;
wire \AXI4Interconnect/_0827_ ;
wire \AXI4Interconnect/_0828_ ;
wire \AXI4Interconnect/_0829_ ;
wire \AXI4Interconnect/_0830_ ;
wire \AXI4Interconnect/_0831_ ;
wire \AXI4Interconnect/_0832_ ;
wire \AXI4Interconnect/_0833_ ;
wire \AXI4Interconnect/_0834_ ;
wire \AXI4Interconnect/_0835_ ;
wire \AXI4Interconnect/_0836_ ;
wire \AXI4Interconnect/_0837_ ;
wire \AXI4Interconnect/_0838_ ;
wire \AXI4Interconnect/_0839_ ;
wire \AXI4Interconnect/_0840_ ;
wire \AXI4Interconnect/_0841_ ;
wire \AXI4Interconnect/_0842_ ;
wire \AXI4Interconnect/_0843_ ;
wire \AXI4Interconnect/_0844_ ;
wire \AXI4Interconnect/_0845_ ;
wire \AXI4Interconnect/_0846_ ;
wire \AXI4Interconnect/_0847_ ;
wire \AXI4Interconnect/_0848_ ;
wire \AXI4Interconnect/_0849_ ;
wire \AXI4Interconnect/_0850_ ;
wire \AXI4Interconnect/_0851_ ;
wire \AXI4Interconnect/_0852_ ;
wire \AXI4Interconnect/_0853_ ;
wire \AXI4Interconnect/_0854_ ;
wire \AXI4Interconnect/_0855_ ;
wire \AXI4Interconnect/_0856_ ;
wire \AXI4Interconnect/_0857_ ;
wire \AXI4Interconnect/_0858_ ;
wire \AXI4Interconnect/_0859_ ;
wire \AXI4Interconnect/_0860_ ;
wire \AXI4Interconnect/_0861_ ;
wire \AXI4Interconnect/_0862_ ;
wire \AXI4Interconnect/_0863_ ;
wire \AXI4Interconnect/_0864_ ;
wire \AXI4Interconnect/_0865_ ;
wire \AXI4Interconnect/_0866_ ;
wire \AXI4Interconnect/_0867_ ;
wire \AXI4Interconnect/_0868_ ;
wire \AXI4Interconnect/_0869_ ;
wire \AXI4Interconnect/_0870_ ;
wire \AXI4Interconnect/_0871_ ;
wire \AXI4Interconnect/_0872_ ;
wire \AXI4Interconnect/_0873_ ;
wire \AXI4Interconnect/_0874_ ;
wire \AXI4Interconnect/_0875_ ;
wire \AXI4Interconnect/_0876_ ;
wire \AXI4Interconnect/_0877_ ;
wire \AXI4Interconnect/_0878_ ;
wire \AXI4Interconnect/_0879_ ;
wire \AXI4Interconnect/_0880_ ;
wire \AXI4Interconnect/_GEN_13 ;
wire \AXI4Interconnect/_GEN_14 ;
wire \AXI4Interconnect/outSelect ;
wire \AXI4Interconnect/selectedReg ;
wire \CLINT/_0000_ ;
wire \CLINT/_0001_ ;
wire \CLINT/_0002_ ;
wire \CLINT/_0003_ ;
wire \CLINT/_0004_ ;
wire \CLINT/_0005_ ;
wire \CLINT/_0006_ ;
wire \CLINT/_0007_ ;
wire \CLINT/_0008_ ;
wire \CLINT/_0009_ ;
wire \CLINT/_0010_ ;
wire \CLINT/_0011_ ;
wire \CLINT/_0012_ ;
wire \CLINT/_0013_ ;
wire \CLINT/_0014_ ;
wire \CLINT/_0015_ ;
wire \CLINT/_0016_ ;
wire \CLINT/_0017_ ;
wire \CLINT/_0018_ ;
wire \CLINT/_0019_ ;
wire \CLINT/_0020_ ;
wire \CLINT/_0021_ ;
wire \CLINT/_0022_ ;
wire \CLINT/_0023_ ;
wire \CLINT/_0024_ ;
wire \CLINT/_0025_ ;
wire \CLINT/_0026_ ;
wire \CLINT/_0027_ ;
wire \CLINT/_0028_ ;
wire \CLINT/_0029_ ;
wire \CLINT/_0030_ ;
wire \CLINT/_0031_ ;
wire \CLINT/_0032_ ;
wire \CLINT/_0033_ ;
wire \CLINT/_0034_ ;
wire \CLINT/_0035_ ;
wire \CLINT/_0036_ ;
wire \CLINT/_0037_ ;
wire \CLINT/_0038_ ;
wire \CLINT/_0039_ ;
wire \CLINT/_0040_ ;
wire \CLINT/_0041_ ;
wire \CLINT/_0042_ ;
wire \CLINT/_0043_ ;
wire \CLINT/_0044_ ;
wire \CLINT/_0045_ ;
wire \CLINT/_0046_ ;
wire \CLINT/_0047_ ;
wire \CLINT/_0048_ ;
wire \CLINT/_0049_ ;
wire \CLINT/_0050_ ;
wire \CLINT/_0051_ ;
wire \CLINT/_0052_ ;
wire \CLINT/_0053_ ;
wire \CLINT/_0054_ ;
wire \CLINT/_0055_ ;
wire \CLINT/_0056_ ;
wire \CLINT/_0057_ ;
wire \CLINT/_0058_ ;
wire \CLINT/_0059_ ;
wire \CLINT/_0060_ ;
wire \CLINT/_0061_ ;
wire \CLINT/_0062_ ;
wire \CLINT/_0063_ ;
wire \CLINT/_0064_ ;
wire \CLINT/_0065_ ;
wire \CLINT/_0066_ ;
wire \CLINT/_0067_ ;
wire \CLINT/_0068_ ;
wire \CLINT/_0069_ ;
wire \CLINT/_0070_ ;
wire \CLINT/_0071_ ;
wire \CLINT/_0072_ ;
wire \CLINT/_0073_ ;
wire \CLINT/_0074_ ;
wire \CLINT/_0075_ ;
wire \CLINT/_0076_ ;
wire \CLINT/_0077_ ;
wire \CLINT/_0078_ ;
wire \CLINT/_0079_ ;
wire \CLINT/_0080_ ;
wire \CLINT/_0081_ ;
wire \CLINT/_0082_ ;
wire \CLINT/_0083_ ;
wire \CLINT/_0084_ ;
wire \CLINT/_0085_ ;
wire \CLINT/_0086_ ;
wire \CLINT/_0087_ ;
wire \CLINT/_0088_ ;
wire \CLINT/_0089_ ;
wire \CLINT/_0090_ ;
wire \CLINT/_0091_ ;
wire \CLINT/_0092_ ;
wire \CLINT/_0093_ ;
wire \CLINT/_0094_ ;
wire \CLINT/_0095_ ;
wire \CLINT/_0096_ ;
wire \CLINT/_0097_ ;
wire \CLINT/_0098_ ;
wire \CLINT/_0099_ ;
wire \CLINT/_0100_ ;
wire \CLINT/_0101_ ;
wire \CLINT/_0102_ ;
wire \CLINT/_0103_ ;
wire \CLINT/_0104_ ;
wire \CLINT/_0105_ ;
wire \CLINT/_0106_ ;
wire \CLINT/_0107_ ;
wire \CLINT/_0108_ ;
wire \CLINT/_0109_ ;
wire \CLINT/_0110_ ;
wire \CLINT/_0111_ ;
wire \CLINT/_0112_ ;
wire \CLINT/_0113_ ;
wire \CLINT/_0114_ ;
wire \CLINT/_0115_ ;
wire \CLINT/_0116_ ;
wire \CLINT/_0117_ ;
wire \CLINT/_0118_ ;
wire \CLINT/_0119_ ;
wire \CLINT/_0120_ ;
wire \CLINT/_0121_ ;
wire \CLINT/_0122_ ;
wire \CLINT/_0123_ ;
wire \CLINT/_0124_ ;
wire \CLINT/_0125_ ;
wire \CLINT/_0126_ ;
wire \CLINT/_0127_ ;
wire \CLINT/_0128_ ;
wire \CLINT/_0129_ ;
wire \CLINT/_0130_ ;
wire \CLINT/_0131_ ;
wire \CLINT/_0132_ ;
wire \CLINT/_0133_ ;
wire \CLINT/_0134_ ;
wire \CLINT/_0135_ ;
wire \CLINT/_0136_ ;
wire \CLINT/_0137_ ;
wire \CLINT/_0138_ ;
wire \CLINT/_0139_ ;
wire \CLINT/_0140_ ;
wire \CLINT/_0141_ ;
wire \CLINT/_0142_ ;
wire \CLINT/_0143_ ;
wire \CLINT/_0144_ ;
wire \CLINT/_0145_ ;
wire \CLINT/_0146_ ;
wire \CLINT/_0147_ ;
wire \CLINT/_0148_ ;
wire \CLINT/_0149_ ;
wire \CLINT/_0150_ ;
wire \CLINT/_0151_ ;
wire \CLINT/_0152_ ;
wire \CLINT/_0153_ ;
wire \CLINT/_0154_ ;
wire \CLINT/_0155_ ;
wire \CLINT/_0156_ ;
wire \CLINT/_0157_ ;
wire \CLINT/_0158_ ;
wire \CLINT/_0159_ ;
wire \CLINT/_0160_ ;
wire \CLINT/_0161_ ;
wire \CLINT/_0162_ ;
wire \CLINT/_0163_ ;
wire \CLINT/_0164_ ;
wire \CLINT/_0165_ ;
wire \CLINT/_0166_ ;
wire \CLINT/_0167_ ;
wire \CLINT/_0168_ ;
wire \CLINT/_0169_ ;
wire \CLINT/_0170_ ;
wire \CLINT/_0171_ ;
wire \CLINT/_0172_ ;
wire \CLINT/_0173_ ;
wire \CLINT/_0174_ ;
wire \CLINT/_0175_ ;
wire \CLINT/_0176_ ;
wire \CLINT/_0177_ ;
wire \CLINT/_0178_ ;
wire \CLINT/_0179_ ;
wire \CLINT/_0180_ ;
wire \CLINT/_0181_ ;
wire \CLINT/_0182_ ;
wire \CLINT/_0183_ ;
wire \CLINT/_0184_ ;
wire \CLINT/_0185_ ;
wire \CLINT/_0186_ ;
wire \CLINT/_0187_ ;
wire \CLINT/_0188_ ;
wire \CLINT/_0189_ ;
wire \CLINT/_0190_ ;
wire \CLINT/_0191_ ;
wire \CLINT/_0192_ ;
wire \CLINT/_0193_ ;
wire \CLINT/_0194_ ;
wire \CLINT/_0195_ ;
wire \CLINT/_0196_ ;
wire \CLINT/_0197_ ;
wire \CLINT/_0198_ ;
wire \CLINT/_0199_ ;
wire \CLINT/_0200_ ;
wire \CLINT/_0201_ ;
wire \CLINT/_0202_ ;
wire \CLINT/_0203_ ;
wire \CLINT/_0204_ ;
wire \CLINT/_0205_ ;
wire \CLINT/_0206_ ;
wire \CLINT/_0207_ ;
wire \CLINT/_0208_ ;
wire \CLINT/_0209_ ;
wire \CLINT/_0210_ ;
wire \CLINT/_0211_ ;
wire \CLINT/_0212_ ;
wire \CLINT/_0213_ ;
wire \CLINT/_0214_ ;
wire \CLINT/_0215_ ;
wire \CLINT/_0216_ ;
wire \CLINT/_0217_ ;
wire \CLINT/_0218_ ;
wire \CLINT/_0219_ ;
wire \CLINT/_0220_ ;
wire \CLINT/_0221_ ;
wire \CLINT/_0222_ ;
wire \CLINT/_0223_ ;
wire \CLINT/_0224_ ;
wire \CLINT/_0225_ ;
wire \CLINT/_0226_ ;
wire \CLINT/_0227_ ;
wire \CLINT/_0228_ ;
wire \CLINT/_0229_ ;
wire \CLINT/_0230_ ;
wire \CLINT/_0231_ ;
wire \CLINT/_0232_ ;
wire \CLINT/_0233_ ;
wire \CLINT/_0234_ ;
wire \CLINT/_0235_ ;
wire \CLINT/_0236_ ;
wire \CLINT/_0237_ ;
wire \CLINT/_0238_ ;
wire \CLINT/_0239_ ;
wire \CLINT/_0240_ ;
wire \CLINT/_0241_ ;
wire \CLINT/_0242_ ;
wire \CLINT/_0243_ ;
wire \CLINT/_0244_ ;
wire \CLINT/_0245_ ;
wire \CLINT/_0246_ ;
wire \CLINT/_0247_ ;
wire \CLINT/_0248_ ;
wire \CLINT/_0249_ ;
wire \CLINT/_0250_ ;
wire \CLINT/_0251_ ;
wire \CLINT/_0252_ ;
wire \CLINT/_0253_ ;
wire \CLINT/_0254_ ;
wire \CLINT/_0255_ ;
wire \CLINT/_0256_ ;
wire \CLINT/_0257_ ;
wire \CLINT/_0258_ ;
wire \CLINT/_0259_ ;
wire \CLINT/_0260_ ;
wire \CLINT/_0261_ ;
wire \CLINT/_0262_ ;
wire \CLINT/_0263_ ;
wire \CLINT/_0264_ ;
wire \CLINT/_0265_ ;
wire \CLINT/_0266_ ;
wire \CLINT/_0267_ ;
wire \CLINT/_0268_ ;
wire \CLINT/_0269_ ;
wire \CLINT/_0270_ ;
wire \CLINT/_0271_ ;
wire \CLINT/_0272_ ;
wire \CLINT/_0273_ ;
wire \CLINT/_0274_ ;
wire \CLINT/_0275_ ;
wire \CLINT/_0276_ ;
wire \CLINT/_0277_ ;
wire \CLINT/_0278_ ;
wire \CLINT/_0279_ ;
wire \CLINT/_0280_ ;
wire \CLINT/_0281_ ;
wire \CLINT/_0282_ ;
wire \CLINT/_0283_ ;
wire \CLINT/_0284_ ;
wire \CLINT/_0285_ ;
wire \CLINT/_0286_ ;
wire \CLINT/_0287_ ;
wire \CLINT/_0288_ ;
wire \CLINT/_0289_ ;
wire \CLINT/_0290_ ;
wire \CLINT/_0291_ ;
wire \CLINT/_0292_ ;
wire \CLINT/_0293_ ;
wire \CLINT/_0294_ ;
wire \CLINT/_0295_ ;
wire \CLINT/_0296_ ;
wire \CLINT/_0297_ ;
wire \CLINT/_0298_ ;
wire \CLINT/_0299_ ;
wire \CLINT/_0300_ ;
wire \CLINT/_0301_ ;
wire \CLINT/_0302_ ;
wire \CLINT/_0303_ ;
wire \CLINT/_0304_ ;
wire \CLINT/_0305_ ;
wire \CLINT/_0306_ ;
wire \CLINT/_0307_ ;
wire \CLINT/_0308_ ;
wire \CLINT/_0309_ ;
wire \CLINT/_0310_ ;
wire \CLINT/_0311_ ;
wire \CLINT/_0312_ ;
wire \CLINT/_0313_ ;
wire \CLINT/_0314_ ;
wire \CLINT/_0315_ ;
wire \CLINT/_0316_ ;
wire \CLINT/_0317_ ;
wire \CLINT/_0318_ ;
wire \CLINT/_0319_ ;
wire \CLINT/_0320_ ;
wire \CLINT/_0321_ ;
wire \CLINT/_0322_ ;
wire \CLINT/_0323_ ;
wire \CLINT/_0324_ ;
wire \CLINT/_0325_ ;
wire \CLINT/_0326_ ;
wire \CLINT/_0327_ ;
wire \CLINT/_0328_ ;
wire \CLINT/_0329_ ;
wire \CLINT/_0330_ ;
wire \CLINT/_0331_ ;
wire \CLINT/_0332_ ;
wire \CLINT/_0333_ ;
wire \CLINT/_0334_ ;
wire \CLINT/_0335_ ;
wire \CLINT/_0336_ ;
wire \CLINT/_0337_ ;
wire \CLINT/_0338_ ;
wire \CLINT/_0339_ ;
wire \CLINT/_0340_ ;
wire \CLINT/_0341_ ;
wire \CLINT/_0342_ ;
wire \CLINT/_0343_ ;
wire \CLINT/_0344_ ;
wire \CLINT/_0345_ ;
wire \CLINT/_0346_ ;
wire \CLINT/_0347_ ;
wire \CLINT/_0348_ ;
wire \CLINT/_0349_ ;
wire \CLINT/_0350_ ;
wire \CLINT/_0351_ ;
wire \CLINT/_0352_ ;
wire \CLINT/_0353_ ;
wire \CLINT/_0354_ ;
wire \CLINT/_0355_ ;
wire \CLINT/_0356_ ;
wire \CLINT/_0357_ ;
wire \CLINT/_0358_ ;
wire \CLINT/_0359_ ;
wire \CLINT/_0360_ ;
wire \CLINT/_0361_ ;
wire \CLINT/_0362_ ;
wire \CLINT/_0363_ ;
wire \CLINT/_0364_ ;
wire \CLINT/_0365_ ;
wire \CLINT/_0366_ ;
wire \CLINT/_0367_ ;
wire \CLINT/_0368_ ;
wire \CLINT/_0369_ ;
wire \CLINT/_0370_ ;
wire \CLINT/_0371_ ;
wire \CLINT/_0372_ ;
wire \CLINT/_0373_ ;
wire \CLINT/_0374_ ;
wire \CLINT/_0375_ ;
wire \CLINT/_0376_ ;
wire \CLINT/_0377_ ;
wire \CLINT/_0378_ ;
wire \CLINT/_0379_ ;
wire \CLINT/_0380_ ;
wire \CLINT/_0381_ ;
wire \CLINT/_0382_ ;
wire \CLINT/_0383_ ;
wire \CLINT/_0384_ ;
wire \CLINT/_0385_ ;
wire \CLINT/_0386_ ;
wire \CLINT/_0387_ ;
wire \CLINT/_0388_ ;
wire \CLINT/_0389_ ;
wire \CLINT/_0390_ ;
wire \CLINT/_0391_ ;
wire \CLINT/_0392_ ;
wire \CLINT/_0393_ ;
wire \CLINT/_0394_ ;
wire \CLINT/_0395_ ;
wire \CLINT/_0396_ ;
wire \CLINT/_0397_ ;
wire \CLINT/_0398_ ;
wire \CLINT/_0399_ ;
wire \CLINT/_0400_ ;
wire \CLINT/_0401_ ;
wire \CLINT/_0402_ ;
wire \CLINT/_0403_ ;
wire \CLINT/_0404_ ;
wire \CLINT/_0405_ ;
wire \CLINT/_0406_ ;
wire \CLINT/_0407_ ;
wire \CLINT/_0408_ ;
wire \CLINT/_0409_ ;
wire \CLINT/_0410_ ;
wire \CLINT/_0411_ ;
wire \CLINT/_0412_ ;
wire \CLINT/_0413_ ;
wire \CLINT/_0414_ ;
wire \CLINT/_0415_ ;
wire \CLINT/_0416_ ;
wire \CLINT/_0417_ ;
wire \CLINT/_0418_ ;
wire \CLINT/_0419_ ;
wire \CLINT/_0420_ ;
wire \CLINT/_0421_ ;
wire \CLINT/_0422_ ;
wire \CLINT/_0423_ ;
wire \CLINT/_0424_ ;
wire \CLINT/_0425_ ;
wire \CLINT/_0426_ ;
wire \CLINT/_0427_ ;
wire \CLINT/_0428_ ;
wire \CLINT/_0429_ ;
wire \CLINT/_0430_ ;
wire \CLINT/_0431_ ;
wire \CLINT/_0432_ ;
wire \CLINT/_0433_ ;
wire \CLINT/_0434_ ;
wire \CLINT/_0435_ ;
wire \CLINT/_0436_ ;
wire \CLINT/_0437_ ;
wire \CLINT/_0438_ ;
wire \CLINT/_0439_ ;
wire \CLINT/_0440_ ;
wire \CLINT/_0441_ ;
wire \CLINT/_0442_ ;
wire \CLINT/_0443_ ;
wire \CLINT/_0444_ ;
wire \CLINT/_0445_ ;
wire \CLINT/_0446_ ;
wire \CLINT/_0447_ ;
wire \CLINT/_0448_ ;
wire \CLINT/_0449_ ;
wire \CLINT/_0450_ ;
wire \CLINT/_0451_ ;
wire \CLINT/_0452_ ;
wire \CLINT/_0453_ ;
wire \CLINT/_0454_ ;
wire \CLINT/_0455_ ;
wire \CLINT/_0456_ ;
wire \CLINT/_0457_ ;
wire \CLINT/_0458_ ;
wire \CLINT/_0459_ ;
wire \CLINT/_0460_ ;
wire \CLINT/_0461_ ;
wire \CLINT/_0462_ ;
wire \CLINT/_0463_ ;
wire \CLINT/_0464_ ;
wire \CLINT/_0465_ ;
wire \CLINT/_0466_ ;
wire \CLINT/_0467_ ;
wire \CLINT/_0468_ ;
wire \CLINT/_0469_ ;
wire \CLINT/_0470_ ;
wire \CLINT/_0471_ ;
wire \CLINT/_0472_ ;
wire \CLINT/_0473_ ;
wire \CLINT/_0474_ ;
wire \CLINT/_0475_ ;
wire \CLINT/_0476_ ;
wire \CLINT/_0477_ ;
wire \CLINT/_0478_ ;
wire \CLINT/_0479_ ;
wire \CLINT/_0480_ ;
wire \CLINT/_0481_ ;
wire \CLINT/_0482_ ;
wire \CLINT/_0483_ ;
wire \CLINT/_0484_ ;
wire \CLINT/_0485_ ;
wire \CLINT/_0486_ ;
wire \CLINT/_0487_ ;
wire \CLINT/_0488_ ;
wire \CLINT/_0489_ ;
wire \CLINT/_0490_ ;
wire \CLINT/_0491_ ;
wire \CLINT/_0492_ ;
wire \CLINT/_0493_ ;
wire \CLINT/_0494_ ;
wire \CLINT/_0495_ ;
wire \CLINT/_0496_ ;
wire \CLINT/_0497_ ;
wire \CLINT/_0498_ ;
wire \CLINT/_0499_ ;
wire \CLINT/_0500_ ;
wire \CLINT/_0501_ ;
wire \CLINT/_0502_ ;
wire \CLINT/_0503_ ;
wire \CLINT/_0504_ ;
wire \CLINT/_0505_ ;
wire \CLINT/_0506_ ;
wire \CLINT/_0507_ ;
wire \CLINT/_0508_ ;
wire \CLINT/_0509_ ;
wire \CLINT/_0510_ ;
wire \CLINT/_0511_ ;
wire \CLINT/_0512_ ;
wire \CLINT/_0513_ ;
wire \CLINT/_0514_ ;
wire \CLINT/_0515_ ;
wire \CLINT/_0516_ ;
wire \CLINT/_0517_ ;
wire \CLINT/_0518_ ;
wire \CLINT/_0519_ ;
wire \CLINT/_0520_ ;
wire \CLINT/_0521_ ;
wire \CLINT/_0522_ ;
wire \CLINT/_0523_ ;
wire \CLINT/_0524_ ;
wire \CLINT/_0525_ ;
wire \CLINT/_0526_ ;
wire \CLINT/_0527_ ;
wire \CLINT/_0528_ ;
wire \CLINT/_0529_ ;
wire \CLINT/_0530_ ;
wire \CLINT/_0531_ ;
wire \CLINT/_0532_ ;
wire \CLINT/_0533_ ;
wire \CLINT/_0534_ ;
wire \CLINT/_0535_ ;
wire \CLINT/_0536_ ;
wire \CLINT/_0537_ ;
wire \CLINT/_0538_ ;
wire \CLINT/_0539_ ;
wire \CLINT/_0540_ ;
wire \CLINT/_0541_ ;
wire \CLINT/_0542_ ;
wire \CLINT/_0543_ ;
wire \CLINT/_0544_ ;
wire \CLINT/_0545_ ;
wire \CLINT/_0546_ ;
wire \CLINT/_0547_ ;
wire \CLINT/_0548_ ;
wire \CLINT/_0549_ ;
wire \CLINT/_0550_ ;
wire \CLINT/_0551_ ;
wire \CLINT/_0552_ ;
wire \CLINT/_0553_ ;
wire \CLINT/_0554_ ;
wire \CLINT/_0555_ ;
wire \CLINT/_0556_ ;
wire \CLINT/_0557_ ;
wire \CLINT/_0558_ ;
wire \CLINT/_0559_ ;
wire \CLINT/_0560_ ;
wire \CLINT/_0561_ ;
wire \CLINT/_0562_ ;
wire \CLINT/_0563_ ;
wire \CLINT/_0564_ ;
wire \CLINT/_0565_ ;
wire \CLINT/_0566_ ;
wire \CLINT/_0567_ ;
wire \CLINT/_0568_ ;
wire \CLINT/_0569_ ;
wire \CLINT/_0570_ ;
wire \CLINT/_0571_ ;
wire \CLINT/_0572_ ;
wire \CLINT/_0573_ ;
wire \CLINT/_0574_ ;
wire \CLINT/_0575_ ;
wire \CLINT/_0576_ ;
wire \CLINT/_0577_ ;
wire \CLINT/_0578_ ;
wire \CLINT/_0579_ ;
wire \CLINT/_0580_ ;
wire \CLINT/_0581_ ;
wire \CLINT/_0582_ ;
wire \CLINT/_0583_ ;
wire \CLINT/_0584_ ;
wire \CLINT/_0585_ ;
wire \CLINT/_0586_ ;
wire \CLINT/_0587_ ;
wire \CLINT/_0588_ ;
wire \CLINT/_0589_ ;
wire \CLINT/_0590_ ;
wire \CLINT/_0591_ ;
wire \CLINT/_0592_ ;
wire \CLINT/_0593_ ;
wire \CLINT/_0594_ ;
wire \CLINT/_0595_ ;
wire \CLINT/_0596_ ;
wire \CLINT/_0597_ ;
wire \CLINT/_0598_ ;
wire \CLINT/_0599_ ;
wire \CLINT/_0600_ ;
wire \CLINT/_0601_ ;
wire \CLINT/_0602_ ;
wire \CLINT/_0603_ ;
wire \CLINT/_0604_ ;
wire \CLINT/_0605_ ;
wire \CLINT/_0606_ ;
wire \CLINT/_0607_ ;
wire \CLINT/_0608_ ;
wire \CLINT/_0609_ ;
wire \CLINT/_0610_ ;
wire \CLINT/_0611_ ;
wire \CLINT/_0612_ ;
wire \CLINT/_0613_ ;
wire \CLINT/_0614_ ;
wire \CLINT/_0615_ ;
wire \CLINT/_0616_ ;
wire \CLINT/_0617_ ;
wire \CLINT/_0618_ ;
wire \CLINT/_0619_ ;
wire \CLINT/_0620_ ;
wire \CLINT/_0621_ ;
wire \CLINT/_0622_ ;
wire \CLINT/_0623_ ;
wire \CLINT/_0624_ ;
wire \CLINT/_0625_ ;
wire \CLINT/_0626_ ;
wire \CLINT/_0627_ ;
wire \CLINT/_0628_ ;
wire \CLINT/_0629_ ;
wire \CLINT/_0630_ ;
wire \CLINT/_0631_ ;
wire \CLINT/_0632_ ;
wire \CLINT/_0633_ ;
wire \CLINT/_0634_ ;
wire \CLINT/_0635_ ;
wire \CLINT/_0636_ ;
wire \CLINT/_0637_ ;
wire \CLINT/_0638_ ;
wire \CLINT/_0639_ ;
wire \CLINT/_0640_ ;
wire \CLINT/_0641_ ;
wire \CLINT/_0642_ ;
wire \CLINT/_0643_ ;
wire \CLINT/_0644_ ;
wire \CLINT/_0645_ ;
wire \CLINT/_0646_ ;
wire \CLINT/_0647_ ;
wire \CLINT/_0648_ ;
wire \CLINT/_0649_ ;
wire \CLINT/_0650_ ;
wire \CLINT/_0651_ ;
wire \CLINT/_0652_ ;
wire \CLINT/_0653_ ;
wire \CLINT/_0654_ ;
wire \CLINT/_0655_ ;
wire \CLINT/_0656_ ;
wire \CLINT/_0657_ ;
wire \CLINT/_0658_ ;
wire \CLINT/_0659_ ;
wire \CLINT/_0660_ ;
wire \CLINT/_0661_ ;
wire \CLINT/_0662_ ;
wire \CLINT/_0663_ ;
wire \CLINT/_0664_ ;
wire \CLINT/_0665_ ;
wire \CLINT/_0666_ ;
wire \CLINT/_0667_ ;
wire \CLINT/_0668_ ;
wire \CLINT/_0669_ ;
wire \CLINT/_0670_ ;
wire \CLINT/_0671_ ;
wire \CLINT/_0672_ ;
wire \CLINT/_0673_ ;
wire \CLINT/_0674_ ;
wire \CLINT/_0675_ ;
wire \CLINT/_0676_ ;
wire \CLINT/_0677_ ;
wire \CLINT/_0678_ ;
wire \CLINT/_0679_ ;
wire \CLINT/_0680_ ;
wire \CLINT/_0681_ ;
wire \CLINT/_0682_ ;
wire \CLINT/_0683_ ;
wire \CLINT/_0684_ ;
wire \CLINT/_0685_ ;
wire \CLINT/_0686_ ;
wire \CLINT/_0687_ ;
wire \CLINT/_0688_ ;
wire \CLINT/_0689_ ;
wire \CLINT/_0690_ ;
wire \CLINT/_0691_ ;
wire \CLINT/_0692_ ;
wire \CLINT/_0693_ ;
wire \CLINT/_0694_ ;
wire \CLINT/_0695_ ;
wire \CLINT/_0696_ ;
wire \CLINT/_0697_ ;
wire \CLINT/_0698_ ;
wire \CLINT/_0699_ ;
wire \CLINT/_0700_ ;
wire \CLINT/_0701_ ;
wire \CLINT/_0702_ ;
wire \CLINT/_0703_ ;
wire \CLINT/_0704_ ;
wire \CLINT/_0705_ ;
wire \CLINT/_0706_ ;
wire \CLINT/_0707_ ;
wire \CLINT/_0708_ ;
wire \CLINT/_0709_ ;
wire \CLINT/_0710_ ;
wire \CLINT/_0711_ ;
wire \CLINT/_0712_ ;
wire \CLINT/_0713_ ;
wire \CLINT/_0714_ ;
wire \CLINT/_0715_ ;
wire \CLINT/_0716_ ;
wire \CLINT/_0717_ ;
wire \CLINT/_0718_ ;
wire \CLINT/_0719_ ;
wire \CLINT/_0720_ ;
wire \CLINT/_0721_ ;
wire \CLINT/_0722_ ;
wire \CLINT/_0723_ ;
wire \CLINT/_0724_ ;
wire \CLINT/_0725_ ;
wire \CLINT/_0726_ ;
wire \CLINT/_0727_ ;
wire \CLINT/_0728_ ;
wire \CLINT/_0729_ ;
wire \CLINT/_0730_ ;
wire \CLINT/_0731_ ;
wire \CLINT/_0732_ ;
wire \CLINT/_0733_ ;
wire \CLINT/_0734_ ;
wire \CLINT/_0735_ ;
wire \CLINT/_0736_ ;
wire \CLINT/_0737_ ;
wire \CLINT/_0738_ ;
wire \CLINT/_0739_ ;
wire \CLINT/_0740_ ;
wire \CLINT/_0741_ ;
wire \CLINT/_0742_ ;
wire \CLINT/_0743_ ;
wire \CLINT/_0744_ ;
wire \CLINT/_0745_ ;
wire \CLINT/_0746_ ;
wire \CLINT/_0747_ ;
wire \CLINT/_0748_ ;
wire \CLINT/_0749_ ;
wire \CLINT/_0750_ ;
wire \CLINT/_0751_ ;
wire \CLINT/_0752_ ;
wire \CLINT/_0753_ ;
wire \CLINT/_0754_ ;
wire \CLINT/_0755_ ;
wire \CLINT/_0756_ ;
wire \CLINT/_0757_ ;
wire \CLINT/_0758_ ;
wire \CLINT/_0759_ ;
wire \CLINT/_0760_ ;
wire \CLINT/_0761_ ;
wire \CLINT/_0762_ ;
wire \CLINT/_0763_ ;
wire \CLINT/_0764_ ;
wire \CLINT/_0765_ ;
wire \CLINT/_0766_ ;
wire \CLINT/_0767_ ;
wire \CLINT/_0768_ ;
wire \CLINT/_0769_ ;
wire \CLINT/_0770_ ;
wire \CLINT/_0771_ ;
wire \CLINT/_0772_ ;
wire \CLINT/_0773_ ;
wire \CLINT/_0774_ ;
wire \CLINT/_0775_ ;
wire \CLINT/_0776_ ;
wire \CLINT/_0777_ ;
wire \CLINT/_0778_ ;
wire \CLINT/_0779_ ;
wire \CLINT/_0780_ ;
wire \CLINT/_0781_ ;
wire \CLINT/_0782_ ;
wire \CLINT/_0783_ ;
wire \CLINT/_0784_ ;
wire \CLINT/_0785_ ;
wire \CLINT/_0786_ ;
wire \CLINT/_0787_ ;
wire \CLINT/_0788_ ;
wire \CLINT/_0789_ ;
wire \CLINT/_0790_ ;
wire \CLINT/_0791_ ;
wire \CLINT/_0792_ ;
wire \CLINT/_0793_ ;
wire \CLINT/_0794_ ;
wire \CLINT/_0795_ ;
wire \CLINT/_0796_ ;
wire \CLINT/_0797_ ;
wire \CLINT/_0798_ ;
wire \CLINT/_0799_ ;
wire \CLINT/_0800_ ;
wire \CLINT/_0801_ ;
wire \CLINT/_0802_ ;
wire \CLINT/_0803_ ;
wire \CLINT/_0804_ ;
wire \CLINT/_0805_ ;
wire \CLINT/_0806_ ;
wire \CLINT/_0807_ ;
wire \CLINT/_0808_ ;
wire \CLINT/_0809_ ;
wire \CLINT/_0810_ ;
wire \CLINT/_0811_ ;
wire \CLINT/_0812_ ;
wire \CLINT/_0813_ ;
wire \CLINT/_0814_ ;
wire \CLINT/_0815_ ;
wire \CLINT/_0816_ ;
wire \CLINT/_0817_ ;
wire \CLINT/_0818_ ;
wire \CLINT/_0819_ ;
wire \CLINT/_0820_ ;
wire \CLINT/_0821_ ;
wire \CLINT/_0822_ ;
wire \CLINT/_0823_ ;
wire \CLINT/_0824_ ;
wire \CLINT/_0825_ ;
wire \CLINT/_0826_ ;
wire \CLINT/_0827_ ;
wire \CLINT/_0828_ ;
wire \CLINT/_0829_ ;
wire \CLINT/_0830_ ;
wire \CLINT/_0831_ ;
wire \CLINT/_0832_ ;
wire \CLINT/_0833_ ;
wire \CLINT/_0834_ ;
wire \CLINT/_0835_ ;
wire \CLINT/_0836_ ;
wire \CLINT/_0837_ ;
wire \EXU/_0000_ ;
wire \EXU/_0001_ ;
wire \EXU/_0002_ ;
wire \EXU/_0003_ ;
wire \EXU/_0004_ ;
wire \EXU/_0005_ ;
wire \EXU/_0006_ ;
wire \EXU/_0007_ ;
wire \EXU/_0008_ ;
wire \EXU/_0009_ ;
wire \EXU/_0010_ ;
wire \EXU/_0011_ ;
wire \EXU/_0012_ ;
wire \EXU/_0013_ ;
wire \EXU/_0014_ ;
wire \EXU/_0015_ ;
wire \EXU/_0016_ ;
wire \EXU/_0017_ ;
wire \EXU/_0018_ ;
wire \EXU/_0019_ ;
wire \EXU/_0020_ ;
wire \EXU/_0021_ ;
wire \EXU/_0022_ ;
wire \EXU/_0023_ ;
wire \EXU/_0024_ ;
wire \EXU/_0025_ ;
wire \EXU/_0026_ ;
wire \EXU/_0027_ ;
wire \EXU/_0028_ ;
wire \EXU/_0029_ ;
wire \EXU/_0030_ ;
wire \EXU/_0031_ ;
wire \EXU/_0032_ ;
wire \EXU/_0033_ ;
wire \EXU/_0034_ ;
wire \EXU/_0035_ ;
wire \EXU/_0036_ ;
wire \EXU/_0037_ ;
wire \EXU/_0038_ ;
wire \EXU/_0039_ ;
wire \EXU/_0040_ ;
wire \EXU/_0041_ ;
wire \EXU/_0042_ ;
wire \EXU/_0043_ ;
wire \EXU/_0044_ ;
wire \EXU/_0045_ ;
wire \EXU/_0046_ ;
wire \EXU/_0047_ ;
wire \EXU/_0048_ ;
wire \EXU/_0049_ ;
wire \EXU/_0050_ ;
wire \EXU/_0051_ ;
wire \EXU/_0052_ ;
wire \EXU/_0053_ ;
wire \EXU/_0054_ ;
wire \EXU/_0055_ ;
wire \EXU/_0056_ ;
wire \EXU/_0057_ ;
wire \EXU/_0058_ ;
wire \EXU/_0059_ ;
wire \EXU/_0060_ ;
wire \EXU/_0061_ ;
wire \EXU/_0062_ ;
wire \EXU/_0063_ ;
wire \EXU/_0064_ ;
wire \EXU/_0065_ ;
wire \EXU/_0066_ ;
wire \EXU/_0067_ ;
wire \EXU/_0068_ ;
wire \EXU/_0069_ ;
wire \EXU/_0070_ ;
wire \EXU/_0071_ ;
wire \EXU/_0072_ ;
wire \EXU/_0073_ ;
wire \EXU/_0074_ ;
wire \EXU/_0075_ ;
wire \EXU/_0076_ ;
wire \EXU/_0077_ ;
wire \EXU/_0078_ ;
wire \EXU/_0079_ ;
wire \EXU/_0080_ ;
wire \EXU/_0081_ ;
wire \EXU/_0082_ ;
wire \EXU/_0083_ ;
wire \EXU/_0084_ ;
wire \EXU/_0085_ ;
wire \EXU/_0086_ ;
wire \EXU/_0087_ ;
wire \EXU/_0088_ ;
wire \EXU/_0089_ ;
wire \EXU/_0090_ ;
wire \EXU/_0091_ ;
wire \EXU/_0092_ ;
wire \EXU/_0093_ ;
wire \EXU/_0094_ ;
wire \EXU/_0095_ ;
wire \EXU/_0096_ ;
wire \EXU/_0097_ ;
wire \EXU/_0098_ ;
wire \EXU/_0099_ ;
wire \EXU/_0100_ ;
wire \EXU/_0101_ ;
wire \EXU/_0102_ ;
wire \EXU/_0103_ ;
wire \EXU/_0104_ ;
wire \EXU/_0105_ ;
wire \EXU/_0106_ ;
wire \EXU/_0107_ ;
wire \EXU/_0108_ ;
wire \EXU/_0109_ ;
wire \EXU/_0110_ ;
wire \EXU/_0111_ ;
wire \EXU/_0112_ ;
wire \EXU/_0113_ ;
wire \EXU/_0114_ ;
wire \EXU/_0115_ ;
wire \EXU/_0116_ ;
wire \EXU/_0117_ ;
wire \EXU/_0118_ ;
wire \EXU/_0119_ ;
wire \EXU/_0120_ ;
wire \EXU/_0121_ ;
wire \EXU/_0122_ ;
wire \EXU/_0123_ ;
wire \EXU/_0124_ ;
wire \EXU/_0125_ ;
wire \EXU/_0126_ ;
wire \EXU/_0127_ ;
wire \EXU/_0128_ ;
wire \EXU/_0129_ ;
wire \EXU/_0130_ ;
wire \EXU/_0131_ ;
wire \EXU/_0132_ ;
wire \EXU/_0133_ ;
wire \EXU/_0134_ ;
wire \EXU/_0135_ ;
wire \EXU/_0136_ ;
wire \EXU/_0137_ ;
wire \EXU/_0138_ ;
wire \EXU/_0139_ ;
wire \EXU/_0140_ ;
wire \EXU/_0141_ ;
wire \EXU/_0142_ ;
wire \EXU/_0143_ ;
wire \EXU/_0144_ ;
wire \EXU/_0145_ ;
wire \EXU/_0146_ ;
wire \EXU/_0147_ ;
wire \EXU/_0148_ ;
wire \EXU/_0149_ ;
wire \EXU/_0150_ ;
wire \EXU/_0151_ ;
wire \EXU/_0152_ ;
wire \EXU/_0153_ ;
wire \EXU/_0154_ ;
wire \EXU/_0155_ ;
wire \EXU/_0156_ ;
wire \EXU/_0157_ ;
wire \EXU/_0158_ ;
wire \EXU/_0159_ ;
wire \EXU/_0160_ ;
wire \EXU/_0161_ ;
wire \EXU/_0162_ ;
wire \EXU/_0163_ ;
wire \EXU/_0164_ ;
wire \EXU/_0165_ ;
wire \EXU/_0166_ ;
wire \EXU/_0167_ ;
wire \EXU/_0168_ ;
wire \EXU/_0169_ ;
wire \EXU/_0170_ ;
wire \EXU/_0171_ ;
wire \EXU/_0172_ ;
wire \EXU/_0173_ ;
wire \EXU/_0174_ ;
wire \EXU/_0175_ ;
wire \EXU/_0176_ ;
wire \EXU/_0177_ ;
wire \EXU/_0178_ ;
wire \EXU/_0179_ ;
wire \EXU/_0180_ ;
wire \EXU/_0181_ ;
wire \EXU/_0182_ ;
wire \EXU/_0183_ ;
wire \EXU/_0184_ ;
wire \EXU/_0185_ ;
wire \EXU/_0186_ ;
wire \EXU/_0187_ ;
wire \EXU/_0188_ ;
wire \EXU/_0189_ ;
wire \EXU/_0190_ ;
wire \EXU/_0191_ ;
wire \EXU/_0192_ ;
wire \EXU/_0193_ ;
wire \EXU/_0194_ ;
wire \EXU/_0195_ ;
wire \EXU/_0196_ ;
wire \EXU/_0197_ ;
wire \EXU/_0198_ ;
wire \EXU/_0199_ ;
wire \EXU/_0200_ ;
wire \EXU/_0201_ ;
wire \EXU/_0202_ ;
wire \EXU/_0203_ ;
wire \EXU/_0204_ ;
wire \EXU/_0205_ ;
wire \EXU/_0206_ ;
wire \EXU/_0207_ ;
wire \EXU/_0208_ ;
wire \EXU/_0209_ ;
wire \EXU/_0210_ ;
wire \EXU/_0211_ ;
wire \EXU/_0212_ ;
wire \EXU/_0213_ ;
wire \EXU/_0214_ ;
wire \EXU/_0215_ ;
wire \EXU/_0216_ ;
wire \EXU/_0217_ ;
wire \EXU/_0218_ ;
wire \EXU/_0219_ ;
wire \EXU/_0220_ ;
wire \EXU/_0221_ ;
wire \EXU/_0222_ ;
wire \EXU/_0223_ ;
wire \EXU/_0224_ ;
wire \EXU/_0225_ ;
wire \EXU/_0226_ ;
wire \EXU/_0227_ ;
wire \EXU/_0228_ ;
wire \EXU/_0229_ ;
wire \EXU/_0230_ ;
wire \EXU/_0231_ ;
wire \EXU/_0232_ ;
wire \EXU/_0233_ ;
wire \EXU/_0234_ ;
wire \EXU/_0235_ ;
wire \EXU/_0236_ ;
wire \EXU/_0237_ ;
wire \EXU/_0238_ ;
wire \EXU/_0239_ ;
wire \EXU/_0240_ ;
wire \EXU/_0241_ ;
wire \EXU/_0242_ ;
wire \EXU/_0243_ ;
wire \EXU/_0244_ ;
wire \EXU/_0245_ ;
wire \EXU/_0246_ ;
wire \EXU/_0247_ ;
wire \EXU/_0248_ ;
wire \EXU/_0249_ ;
wire \EXU/_0250_ ;
wire \EXU/_0251_ ;
wire \EXU/_0252_ ;
wire \EXU/_0253_ ;
wire \EXU/_0254_ ;
wire \EXU/_0255_ ;
wire \EXU/_0256_ ;
wire \EXU/_0257_ ;
wire \EXU/_0258_ ;
wire \EXU/_0259_ ;
wire \EXU/_0260_ ;
wire \EXU/_0261_ ;
wire \EXU/_0262_ ;
wire \EXU/_0263_ ;
wire \EXU/_0264_ ;
wire \EXU/_0265_ ;
wire \EXU/_0266_ ;
wire \EXU/_0267_ ;
wire \EXU/_0268_ ;
wire \EXU/_0269_ ;
wire \EXU/_0270_ ;
wire \EXU/_0271_ ;
wire \EXU/_0272_ ;
wire \EXU/_0273_ ;
wire \EXU/_0274_ ;
wire \EXU/_0275_ ;
wire \EXU/_0276_ ;
wire \EXU/_0277_ ;
wire \EXU/_0278_ ;
wire \EXU/_0279_ ;
wire \EXU/_0280_ ;
wire \EXU/_0281_ ;
wire \EXU/_0282_ ;
wire \EXU/_0283_ ;
wire \EXU/_0284_ ;
wire \EXU/_0285_ ;
wire \EXU/_0286_ ;
wire \EXU/_0287_ ;
wire \EXU/_0288_ ;
wire \EXU/_0289_ ;
wire \EXU/_0290_ ;
wire \EXU/_0291_ ;
wire \EXU/_0292_ ;
wire \EXU/_0293_ ;
wire \EXU/_0294_ ;
wire \EXU/_0295_ ;
wire \EXU/_0296_ ;
wire \EXU/_0297_ ;
wire \EXU/_0298_ ;
wire \EXU/_0299_ ;
wire \EXU/_0300_ ;
wire \EXU/_0301_ ;
wire \EXU/_0302_ ;
wire \EXU/_0303_ ;
wire \EXU/_0304_ ;
wire \EXU/_0305_ ;
wire \EXU/_0306_ ;
wire \EXU/_0307_ ;
wire \EXU/_0308_ ;
wire \EXU/_0309_ ;
wire \EXU/_0310_ ;
wire \EXU/_0311_ ;
wire \EXU/_0312_ ;
wire \EXU/_0313_ ;
wire \EXU/_0314_ ;
wire \EXU/_0315_ ;
wire \EXU/_0316_ ;
wire \EXU/_0317_ ;
wire \EXU/_0318_ ;
wire \EXU/_0319_ ;
wire \EXU/_0320_ ;
wire \EXU/_0321_ ;
wire \EXU/_0322_ ;
wire \EXU/_0323_ ;
wire \EXU/_0324_ ;
wire \EXU/_0325_ ;
wire \EXU/_0326_ ;
wire \EXU/_0327_ ;
wire \EXU/_0328_ ;
wire \EXU/_0329_ ;
wire \EXU/_0330_ ;
wire \EXU/_0331_ ;
wire \EXU/_0332_ ;
wire \EXU/_0333_ ;
wire \EXU/_0334_ ;
wire \EXU/_0335_ ;
wire \EXU/_0336_ ;
wire \EXU/_0337_ ;
wire \EXU/_0338_ ;
wire \EXU/_0339_ ;
wire \EXU/_0340_ ;
wire \EXU/_0341_ ;
wire \EXU/_0342_ ;
wire \EXU/_0343_ ;
wire \EXU/_0344_ ;
wire \EXU/_0345_ ;
wire \EXU/_0346_ ;
wire \EXU/_0347_ ;
wire \EXU/_0348_ ;
wire \EXU/_0349_ ;
wire \EXU/_0350_ ;
wire \EXU/_0351_ ;
wire \EXU/_0352_ ;
wire \EXU/_0353_ ;
wire \EXU/_0354_ ;
wire \EXU/_0355_ ;
wire \EXU/_0356_ ;
wire \EXU/_0357_ ;
wire \EXU/_0358_ ;
wire \EXU/_0359_ ;
wire \EXU/_0360_ ;
wire \EXU/_0361_ ;
wire \EXU/_0362_ ;
wire \EXU/_0363_ ;
wire \EXU/_0364_ ;
wire \EXU/_0365_ ;
wire \EXU/_0366_ ;
wire \EXU/_0367_ ;
wire \EXU/_0368_ ;
wire \EXU/_0369_ ;
wire \EXU/_0370_ ;
wire \EXU/_0371_ ;
wire \EXU/_0372_ ;
wire \EXU/_0373_ ;
wire \EXU/_0374_ ;
wire \EXU/_0375_ ;
wire \EXU/_0376_ ;
wire \EXU/_0377_ ;
wire \EXU/_0378_ ;
wire \EXU/_0379_ ;
wire \EXU/_0380_ ;
wire \EXU/_0381_ ;
wire \EXU/_0382_ ;
wire \EXU/_0383_ ;
wire \EXU/_0384_ ;
wire \EXU/_0385_ ;
wire \EXU/_0386_ ;
wire \EXU/_0387_ ;
wire \EXU/_0388_ ;
wire \EXU/_0389_ ;
wire \EXU/_0390_ ;
wire \EXU/_0391_ ;
wire \EXU/_0392_ ;
wire \EXU/_0393_ ;
wire \EXU/_0394_ ;
wire \EXU/_0395_ ;
wire \EXU/_0396_ ;
wire \EXU/_0397_ ;
wire \EXU/_0398_ ;
wire \EXU/_0399_ ;
wire \EXU/_0400_ ;
wire \EXU/_0401_ ;
wire \EXU/_0402_ ;
wire \EXU/_0403_ ;
wire \EXU/_0404_ ;
wire \EXU/_0405_ ;
wire \EXU/_0406_ ;
wire \EXU/_0407_ ;
wire \EXU/_0408_ ;
wire \EXU/_0409_ ;
wire \EXU/_0410_ ;
wire \EXU/_0411_ ;
wire \EXU/_0412_ ;
wire \EXU/_0413_ ;
wire \EXU/_0414_ ;
wire \EXU/_0415_ ;
wire \EXU/_0416_ ;
wire \EXU/_0417_ ;
wire \EXU/_0418_ ;
wire \EXU/_0419_ ;
wire \EXU/_0420_ ;
wire \EXU/_0421_ ;
wire \EXU/_0422_ ;
wire \EXU/_0423_ ;
wire \EXU/_0424_ ;
wire \EXU/_0425_ ;
wire \EXU/_0426_ ;
wire \EXU/_0427_ ;
wire \EXU/_0428_ ;
wire \EXU/_0429_ ;
wire \EXU/_0430_ ;
wire \EXU/_0431_ ;
wire \EXU/_0432_ ;
wire \EXU/_0433_ ;
wire \EXU/_0434_ ;
wire \EXU/_0435_ ;
wire \EXU/_0436_ ;
wire \EXU/_0437_ ;
wire \EXU/_0438_ ;
wire \EXU/_0439_ ;
wire \EXU/_0440_ ;
wire \EXU/_0441_ ;
wire \EXU/_0442_ ;
wire \EXU/_0443_ ;
wire \EXU/_0444_ ;
wire \EXU/_0445_ ;
wire \EXU/_0446_ ;
wire \EXU/_0447_ ;
wire \EXU/_0448_ ;
wire \EXU/_0449_ ;
wire \EXU/_0450_ ;
wire \EXU/_0451_ ;
wire \EXU/_0452_ ;
wire \EXU/_0453_ ;
wire \EXU/_0454_ ;
wire \EXU/_0455_ ;
wire \EXU/_0456_ ;
wire \EXU/_0457_ ;
wire \EXU/_0458_ ;
wire \EXU/_0459_ ;
wire \EXU/_0460_ ;
wire \EXU/_0461_ ;
wire \EXU/_0462_ ;
wire \EXU/_0463_ ;
wire \EXU/_0464_ ;
wire \EXU/_0465_ ;
wire \EXU/_0466_ ;
wire \EXU/_0467_ ;
wire \EXU/_0468_ ;
wire \EXU/_0469_ ;
wire \EXU/_0470_ ;
wire \EXU/_0471_ ;
wire \EXU/_0472_ ;
wire \EXU/_0473_ ;
wire \EXU/_0474_ ;
wire \EXU/_0475_ ;
wire \EXU/_0476_ ;
wire \EXU/_0477_ ;
wire \EXU/_0478_ ;
wire \EXU/_0479_ ;
wire \EXU/_0480_ ;
wire \EXU/_0481_ ;
wire \EXU/_0482_ ;
wire \EXU/_0483_ ;
wire \EXU/_0484_ ;
wire \EXU/_0485_ ;
wire \EXU/_0486_ ;
wire \EXU/_0487_ ;
wire \EXU/_0488_ ;
wire \EXU/_0489_ ;
wire \EXU/_0490_ ;
wire \EXU/_0491_ ;
wire \EXU/_0492_ ;
wire \EXU/_0493_ ;
wire \EXU/_0494_ ;
wire \EXU/_0495_ ;
wire \EXU/_0496_ ;
wire \EXU/_0497_ ;
wire \EXU/_0498_ ;
wire \EXU/_0499_ ;
wire \EXU/_0500_ ;
wire \EXU/_0501_ ;
wire \EXU/_0502_ ;
wire \EXU/_0503_ ;
wire \EXU/_0504_ ;
wire \EXU/_0505_ ;
wire \EXU/_0506_ ;
wire \EXU/_0507_ ;
wire \EXU/_0508_ ;
wire \EXU/_0509_ ;
wire \EXU/_0510_ ;
wire \EXU/_0511_ ;
wire \EXU/_0512_ ;
wire \EXU/_0513_ ;
wire \EXU/_0514_ ;
wire \EXU/_0515_ ;
wire \EXU/_0516_ ;
wire \EXU/_0517_ ;
wire \EXU/_0518_ ;
wire \EXU/_0519_ ;
wire \EXU/_0520_ ;
wire \EXU/_0521_ ;
wire \EXU/_0522_ ;
wire \EXU/_0523_ ;
wire \EXU/_0524_ ;
wire \EXU/_0525_ ;
wire \EXU/_0526_ ;
wire \EXU/_0527_ ;
wire \EXU/_0528_ ;
wire \EXU/_0529_ ;
wire \EXU/_0530_ ;
wire \EXU/_0531_ ;
wire \EXU/_0532_ ;
wire \EXU/_0533_ ;
wire \EXU/_0534_ ;
wire \EXU/_0535_ ;
wire \EXU/_0536_ ;
wire \EXU/_0537_ ;
wire \EXU/_0538_ ;
wire \EXU/_0539_ ;
wire \EXU/_0540_ ;
wire \EXU/_0541_ ;
wire \EXU/_0542_ ;
wire \EXU/_0543_ ;
wire \EXU/_0544_ ;
wire \EXU/_0545_ ;
wire \EXU/_0546_ ;
wire \EXU/_0547_ ;
wire \EXU/_0548_ ;
wire \EXU/_0549_ ;
wire \EXU/_0550_ ;
wire \EXU/_0551_ ;
wire \EXU/_0552_ ;
wire \EXU/_0553_ ;
wire \EXU/_0554_ ;
wire \EXU/_0555_ ;
wire \EXU/_0556_ ;
wire \EXU/_0557_ ;
wire \EXU/_0558_ ;
wire \EXU/_0559_ ;
wire \EXU/_0560_ ;
wire \EXU/_0561_ ;
wire \EXU/_0562_ ;
wire \EXU/_0563_ ;
wire \EXU/_0564_ ;
wire \EXU/_0565_ ;
wire \EXU/_0566_ ;
wire \EXU/_0567_ ;
wire \EXU/_0568_ ;
wire \EXU/_0569_ ;
wire \EXU/_0570_ ;
wire \EXU/_0571_ ;
wire \EXU/_0572_ ;
wire \EXU/_0573_ ;
wire \EXU/_0574_ ;
wire \EXU/_0575_ ;
wire \EXU/_0576_ ;
wire \EXU/_0577_ ;
wire \EXU/_0578_ ;
wire \EXU/_0579_ ;
wire \EXU/_0580_ ;
wire \EXU/_0581_ ;
wire \EXU/_0582_ ;
wire \EXU/_0583_ ;
wire \EXU/_0584_ ;
wire \EXU/_0585_ ;
wire \EXU/_0586_ ;
wire \EXU/_0587_ ;
wire \EXU/_0588_ ;
wire \EXU/_0589_ ;
wire \EXU/_0590_ ;
wire \EXU/_0591_ ;
wire \EXU/_0592_ ;
wire \EXU/_0593_ ;
wire \EXU/_0594_ ;
wire \EXU/_0595_ ;
wire \EXU/_0596_ ;
wire \EXU/_0597_ ;
wire \EXU/_0598_ ;
wire \EXU/_0599_ ;
wire \EXU/_0600_ ;
wire \EXU/_0601_ ;
wire \EXU/_0602_ ;
wire \EXU/_0603_ ;
wire \EXU/_0604_ ;
wire \EXU/_0605_ ;
wire \EXU/_0606_ ;
wire \EXU/_0607_ ;
wire \EXU/_0608_ ;
wire \EXU/_0609_ ;
wire \EXU/_0610_ ;
wire \EXU/_0611_ ;
wire \EXU/_0612_ ;
wire \EXU/_0613_ ;
wire \EXU/_0614_ ;
wire \EXU/_0615_ ;
wire \EXU/_0616_ ;
wire \EXU/_0617_ ;
wire \EXU/_0618_ ;
wire \EXU/_0619_ ;
wire \EXU/_0620_ ;
wire \EXU/_0621_ ;
wire \EXU/_0622_ ;
wire \EXU/_0623_ ;
wire \EXU/_0624_ ;
wire \EXU/_0625_ ;
wire \EXU/_0626_ ;
wire \EXU/_0627_ ;
wire \EXU/_0628_ ;
wire \EXU/_0629_ ;
wire \EXU/_0630_ ;
wire \EXU/_0631_ ;
wire \EXU/_0632_ ;
wire \EXU/_0633_ ;
wire \EXU/_0634_ ;
wire \EXU/_0635_ ;
wire \EXU/_0636_ ;
wire \EXU/_0637_ ;
wire \EXU/_0638_ ;
wire \EXU/_0639_ ;
wire \EXU/_0640_ ;
wire \EXU/_0641_ ;
wire \EXU/_0642_ ;
wire \EXU/_0643_ ;
wire \EXU/_0644_ ;
wire \EXU/_0645_ ;
wire \EXU/_0646_ ;
wire \EXU/_0647_ ;
wire \EXU/_0648_ ;
wire \EXU/_0649_ ;
wire \EXU/_0650_ ;
wire \EXU/_0651_ ;
wire \EXU/_0652_ ;
wire \EXU/_0653_ ;
wire \EXU/_0654_ ;
wire \EXU/_0655_ ;
wire \EXU/_0656_ ;
wire \EXU/_0657_ ;
wire \EXU/_0658_ ;
wire \EXU/_0659_ ;
wire \EXU/_0660_ ;
wire \EXU/_0661_ ;
wire \EXU/_0662_ ;
wire \EXU/_0663_ ;
wire \EXU/_0664_ ;
wire \EXU/_0665_ ;
wire \EXU/_0666_ ;
wire \EXU/_0667_ ;
wire \EXU/_0668_ ;
wire \EXU/_0669_ ;
wire \EXU/_0670_ ;
wire \EXU/_0671_ ;
wire \EXU/_0672_ ;
wire \EXU/_0673_ ;
wire \EXU/_0674_ ;
wire \EXU/_0675_ ;
wire \EXU/_0676_ ;
wire \EXU/_0677_ ;
wire \EXU/_0678_ ;
wire \EXU/_0679_ ;
wire \EXU/_0680_ ;
wire \EXU/_0681_ ;
wire \EXU/_0682_ ;
wire \EXU/_0683_ ;
wire \EXU/_0684_ ;
wire \EXU/_0685_ ;
wire \EXU/_0686_ ;
wire \EXU/_0687_ ;
wire \EXU/_0688_ ;
wire \EXU/_0689_ ;
wire \EXU/_0690_ ;
wire \EXU/_0691_ ;
wire \EXU/_0692_ ;
wire \EXU/_0693_ ;
wire \EXU/_0694_ ;
wire \EXU/_0695_ ;
wire \EXU/_0696_ ;
wire \EXU/_0697_ ;
wire \EXU/_0698_ ;
wire \EXU/_0699_ ;
wire \EXU/_0700_ ;
wire \EXU/_0701_ ;
wire \EXU/_0702_ ;
wire \EXU/_0703_ ;
wire \EXU/_0704_ ;
wire \EXU/_0705_ ;
wire \EXU/_0706_ ;
wire \EXU/_0707_ ;
wire \EXU/_0708_ ;
wire \EXU/_0709_ ;
wire \EXU/_0710_ ;
wire \EXU/_0711_ ;
wire \EXU/_0712_ ;
wire \EXU/_0713_ ;
wire \EXU/_0714_ ;
wire \EXU/_0715_ ;
wire \EXU/_0716_ ;
wire \EXU/_0717_ ;
wire \EXU/_0718_ ;
wire \EXU/_0719_ ;
wire \EXU/_0720_ ;
wire \EXU/_0721_ ;
wire \EXU/_0722_ ;
wire \EXU/_0723_ ;
wire \EXU/_0724_ ;
wire \EXU/_0725_ ;
wire \EXU/_0726_ ;
wire \EXU/_0727_ ;
wire \EXU/_0728_ ;
wire \EXU/_0729_ ;
wire \EXU/_0730_ ;
wire \EXU/_0731_ ;
wire \EXU/_0732_ ;
wire \EXU/_0733_ ;
wire \EXU/_0734_ ;
wire \EXU/_0735_ ;
wire \EXU/_0736_ ;
wire \EXU/_0737_ ;
wire \EXU/_0738_ ;
wire \EXU/_0739_ ;
wire \EXU/_0740_ ;
wire \EXU/_0741_ ;
wire \EXU/_0742_ ;
wire \EXU/_0743_ ;
wire \EXU/_0744_ ;
wire \EXU/_0745_ ;
wire \EXU/_0746_ ;
wire \EXU/_0747_ ;
wire \EXU/_0748_ ;
wire \EXU/_0749_ ;
wire \EXU/_0750_ ;
wire \EXU/_0751_ ;
wire \EXU/_0752_ ;
wire \EXU/_0753_ ;
wire \EXU/_0754_ ;
wire \EXU/_0755_ ;
wire \EXU/_0756_ ;
wire \EXU/_0757_ ;
wire \EXU/_0758_ ;
wire \EXU/_0759_ ;
wire \EXU/_0760_ ;
wire \EXU/_0761_ ;
wire \EXU/_0762_ ;
wire \EXU/_0763_ ;
wire \EXU/_0764_ ;
wire \EXU/_0765_ ;
wire \EXU/_0766_ ;
wire \EXU/_0767_ ;
wire \EXU/_0768_ ;
wire \EXU/_0769_ ;
wire \EXU/_0770_ ;
wire \EXU/_0771_ ;
wire \EXU/_0772_ ;
wire \EXU/_0773_ ;
wire \EXU/_0774_ ;
wire \EXU/_0775_ ;
wire \EXU/_0776_ ;
wire \EXU/_0777_ ;
wire \EXU/_0778_ ;
wire \EXU/_0779_ ;
wire \EXU/_0780_ ;
wire \EXU/_0781_ ;
wire \EXU/_0782_ ;
wire \EXU/_0783_ ;
wire \EXU/_0784_ ;
wire \EXU/_0785_ ;
wire \EXU/_0786_ ;
wire \EXU/_0787_ ;
wire \EXU/_0788_ ;
wire \EXU/_0789_ ;
wire \EXU/_0790_ ;
wire \EXU/_0791_ ;
wire \EXU/_0792_ ;
wire \EXU/_0793_ ;
wire \EXU/_0794_ ;
wire \EXU/_0795_ ;
wire \EXU/_0796_ ;
wire \EXU/_0797_ ;
wire \EXU/_0798_ ;
wire \EXU/_0799_ ;
wire \EXU/_0800_ ;
wire \EXU/_0801_ ;
wire \EXU/_0802_ ;
wire \EXU/_0803_ ;
wire \EXU/_0804_ ;
wire \EXU/_0805_ ;
wire \EXU/_0806_ ;
wire \EXU/_0807_ ;
wire \EXU/_0808_ ;
wire \EXU/_0809_ ;
wire \EXU/_0810_ ;
wire \EXU/_0811_ ;
wire \EXU/_0812_ ;
wire \EXU/_0813_ ;
wire \EXU/_0814_ ;
wire \EXU/_0815_ ;
wire \EXU/_0816_ ;
wire \EXU/_0817_ ;
wire \EXU/_0818_ ;
wire \EXU/_0819_ ;
wire \EXU/_0820_ ;
wire \EXU/_0821_ ;
wire \EXU/_0822_ ;
wire \EXU/_0823_ ;
wire \EXU/_0824_ ;
wire \EXU/_0825_ ;
wire \EXU/_0826_ ;
wire \EXU/_0827_ ;
wire \EXU/_0828_ ;
wire \EXU/_0829_ ;
wire \EXU/_0830_ ;
wire \EXU/_0831_ ;
wire \EXU/_0832_ ;
wire \EXU/_0833_ ;
wire \EXU/_0834_ ;
wire \EXU/_0835_ ;
wire \EXU/_0836_ ;
wire \EXU/_0837_ ;
wire \EXU/_0838_ ;
wire \EXU/_0839_ ;
wire \EXU/_0840_ ;
wire \EXU/_0841_ ;
wire \EXU/_0842_ ;
wire \EXU/_0843_ ;
wire \EXU/_0844_ ;
wire \EXU/_0845_ ;
wire \EXU/_0846_ ;
wire \EXU/_0847_ ;
wire \EXU/_0848_ ;
wire \EXU/_0849_ ;
wire \EXU/_0850_ ;
wire \EXU/_0851_ ;
wire \EXU/_0852_ ;
wire \EXU/_0853_ ;
wire \EXU/_0854_ ;
wire \EXU/_0855_ ;
wire \EXU/_0856_ ;
wire \EXU/_0857_ ;
wire \EXU/_0858_ ;
wire \EXU/_0859_ ;
wire \EXU/_0860_ ;
wire \EXU/_0861_ ;
wire \EXU/_0862_ ;
wire \EXU/_0863_ ;
wire \EXU/_0864_ ;
wire \EXU/_0865_ ;
wire \EXU/_0866_ ;
wire \EXU/_0867_ ;
wire \EXU/_0868_ ;
wire \EXU/_0869_ ;
wire \EXU/_0870_ ;
wire \EXU/_0871_ ;
wire \EXU/_0872_ ;
wire \EXU/_0873_ ;
wire \EXU/_0874_ ;
wire \EXU/_0875_ ;
wire \EXU/_0876_ ;
wire \EXU/_0877_ ;
wire \EXU/_0878_ ;
wire \EXU/_0879_ ;
wire \EXU/_0880_ ;
wire \EXU/_0881_ ;
wire \EXU/_0882_ ;
wire \EXU/_0883_ ;
wire \EXU/_0884_ ;
wire \EXU/_0885_ ;
wire \EXU/_0886_ ;
wire \EXU/_0887_ ;
wire \EXU/_0888_ ;
wire \EXU/_0889_ ;
wire \EXU/_0890_ ;
wire \EXU/_0891_ ;
wire \EXU/_0892_ ;
wire \EXU/_0893_ ;
wire \EXU/_0894_ ;
wire \EXU/_0895_ ;
wire \EXU/_0896_ ;
wire \EXU/_0897_ ;
wire \EXU/_0898_ ;
wire \EXU/_0899_ ;
wire \EXU/_0900_ ;
wire \EXU/_0901_ ;
wire \EXU/_0902_ ;
wire \EXU/_0903_ ;
wire \EXU/_0904_ ;
wire \EXU/_0905_ ;
wire \EXU/_0906_ ;
wire \EXU/_0907_ ;
wire \EXU/_0908_ ;
wire \EXU/_0909_ ;
wire \EXU/_0910_ ;
wire \EXU/_0911_ ;
wire \EXU/_0912_ ;
wire \EXU/_0913_ ;
wire \EXU/_0914_ ;
wire \EXU/_0915_ ;
wire \EXU/_0916_ ;
wire \EXU/_0917_ ;
wire \EXU/_0918_ ;
wire \EXU/_0919_ ;
wire \EXU/_0920_ ;
wire \EXU/_0921_ ;
wire \EXU/_0922_ ;
wire \EXU/_0923_ ;
wire \EXU/_0924_ ;
wire \EXU/_0925_ ;
wire \EXU/_0926_ ;
wire \EXU/_0927_ ;
wire \EXU/_0928_ ;
wire \EXU/_0929_ ;
wire \EXU/_0930_ ;
wire \EXU/_0931_ ;
wire \EXU/_0932_ ;
wire \EXU/_0933_ ;
wire \EXU/_0934_ ;
wire \EXU/_0935_ ;
wire \EXU/_0936_ ;
wire \EXU/_0937_ ;
wire \EXU/_0938_ ;
wire \EXU/_0939_ ;
wire \EXU/_0940_ ;
wire \EXU/_0941_ ;
wire \EXU/_0942_ ;
wire \EXU/_0943_ ;
wire \EXU/_0944_ ;
wire \EXU/_0945_ ;
wire \EXU/_0946_ ;
wire \EXU/_0947_ ;
wire \EXU/_0948_ ;
wire \EXU/_0949_ ;
wire \EXU/_0950_ ;
wire \EXU/_0951_ ;
wire \EXU/_0952_ ;
wire \EXU/_0953_ ;
wire \EXU/_0954_ ;
wire \EXU/_0955_ ;
wire \EXU/_0956_ ;
wire \EXU/_0957_ ;
wire \EXU/_0958_ ;
wire \EXU/_0959_ ;
wire \EXU/_0960_ ;
wire \EXU/_0961_ ;
wire \EXU/_0962_ ;
wire \EXU/_0963_ ;
wire \EXU/_0964_ ;
wire \EXU/_0965_ ;
wire \EXU/_0966_ ;
wire \EXU/_0967_ ;
wire \EXU/_0968_ ;
wire \EXU/_0969_ ;
wire \EXU/_0970_ ;
wire \EXU/_0971_ ;
wire \EXU/_0972_ ;
wire \EXU/_0973_ ;
wire \EXU/_0974_ ;
wire \EXU/_0975_ ;
wire \EXU/_0976_ ;
wire \EXU/_0977_ ;
wire \EXU/_0978_ ;
wire \EXU/_0979_ ;
wire \EXU/_0980_ ;
wire \EXU/_0981_ ;
wire \EXU/_0982_ ;
wire \EXU/_0983_ ;
wire \EXU/_0984_ ;
wire \EXU/_0985_ ;
wire \EXU/_0986_ ;
wire \EXU/_0987_ ;
wire \EXU/_0988_ ;
wire \EXU/_0989_ ;
wire \EXU/_0990_ ;
wire \EXU/_0991_ ;
wire \EXU/_0992_ ;
wire \EXU/_0993_ ;
wire \EXU/_0994_ ;
wire \EXU/_0995_ ;
wire \EXU/_0996_ ;
wire \EXU/_0997_ ;
wire \EXU/_0998_ ;
wire \EXU/_0999_ ;
wire \EXU/_1000_ ;
wire \EXU/_1001_ ;
wire \EXU/_1002_ ;
wire \EXU/_1003_ ;
wire \EXU/_1004_ ;
wire \EXU/_1005_ ;
wire \EXU/_1006_ ;
wire \EXU/_1007_ ;
wire \EXU/_1008_ ;
wire \EXU/_1009_ ;
wire \EXU/_1010_ ;
wire \EXU/_1011_ ;
wire \EXU/_1012_ ;
wire \EXU/_1013_ ;
wire \EXU/_1014_ ;
wire \EXU/_1015_ ;
wire \EXU/_1016_ ;
wire \EXU/_1017_ ;
wire \EXU/_1018_ ;
wire \EXU/_1019_ ;
wire \EXU/_1020_ ;
wire \EXU/_1021_ ;
wire \EXU/_1022_ ;
wire \EXU/_1023_ ;
wire \EXU/_1024_ ;
wire \EXU/_1025_ ;
wire \EXU/_1026_ ;
wire \EXU/_1027_ ;
wire \EXU/_1028_ ;
wire \EXU/_1029_ ;
wire \EXU/_1030_ ;
wire \EXU/_1031_ ;
wire \EXU/_1032_ ;
wire \EXU/_1033_ ;
wire \EXU/_1034_ ;
wire \EXU/_1035_ ;
wire \EXU/_1036_ ;
wire \EXU/_1037_ ;
wire \EXU/_1038_ ;
wire \EXU/_1039_ ;
wire \EXU/_1040_ ;
wire \EXU/_1041_ ;
wire \EXU/_1042_ ;
wire \EXU/_1043_ ;
wire \EXU/_1044_ ;
wire \EXU/_1045_ ;
wire \EXU/_1046_ ;
wire \EXU/_1047_ ;
wire \EXU/_1048_ ;
wire \EXU/_1049_ ;
wire \EXU/_1050_ ;
wire \EXU/_1051_ ;
wire \EXU/_1052_ ;
wire \EXU/_1053_ ;
wire \EXU/_1054_ ;
wire \EXU/_1055_ ;
wire \EXU/_1056_ ;
wire \EXU/_1057_ ;
wire \EXU/_1058_ ;
wire \EXU/_1059_ ;
wire \EXU/_1060_ ;
wire \EXU/_1061_ ;
wire \EXU/_1062_ ;
wire \EXU/_1063_ ;
wire \EXU/_1064_ ;
wire \EXU/_1065_ ;
wire \EXU/_1066_ ;
wire \EXU/_1067_ ;
wire \EXU/_1068_ ;
wire \EXU/_1069_ ;
wire \EXU/_1070_ ;
wire \EXU/_1071_ ;
wire \EXU/_1072_ ;
wire \EXU/_1073_ ;
wire \EXU/_1074_ ;
wire \EXU/_1075_ ;
wire \EXU/_1076_ ;
wire \EXU/_1077_ ;
wire \EXU/_1078_ ;
wire \EXU/_1079_ ;
wire \EXU/_1080_ ;
wire \EXU/_1081_ ;
wire \EXU/_1082_ ;
wire \EXU/_1083_ ;
wire \EXU/_1084_ ;
wire \EXU/_1085_ ;
wire \EXU/_1086_ ;
wire \EXU/_1087_ ;
wire \EXU/_1088_ ;
wire \EXU/_1089_ ;
wire \EXU/_1090_ ;
wire \EXU/_1091_ ;
wire \EXU/_1092_ ;
wire \EXU/_1093_ ;
wire \EXU/_1094_ ;
wire \EXU/_1095_ ;
wire \EXU/_1096_ ;
wire \EXU/_1097_ ;
wire \EXU/_1098_ ;
wire \EXU/_1099_ ;
wire \EXU/_1100_ ;
wire \EXU/_1101_ ;
wire \EXU/_1102_ ;
wire \EXU/_1103_ ;
wire \EXU/_1104_ ;
wire \EXU/_1105_ ;
wire \EXU/_1106_ ;
wire \EXU/_1107_ ;
wire \EXU/_1108_ ;
wire \EXU/_1109_ ;
wire \EXU/_1110_ ;
wire \EXU/_1111_ ;
wire \EXU/_1112_ ;
wire \EXU/_1113_ ;
wire \EXU/_1114_ ;
wire \EXU/_1115_ ;
wire \EXU/_1116_ ;
wire \EXU/_1117_ ;
wire \EXU/_1118_ ;
wire \EXU/_1119_ ;
wire \EXU/_1120_ ;
wire \EXU/_1121_ ;
wire \EXU/_1122_ ;
wire \EXU/_1123_ ;
wire \EXU/_1124_ ;
wire \EXU/_1125_ ;
wire \EXU/_1126_ ;
wire \EXU/_1127_ ;
wire \EXU/_1128_ ;
wire \EXU/_1129_ ;
wire \EXU/_1130_ ;
wire \EXU/_1131_ ;
wire \EXU/_1132_ ;
wire \EXU/_1133_ ;
wire \EXU/_1134_ ;
wire \EXU/_1135_ ;
wire \EXU/_1136_ ;
wire \EXU/_1137_ ;
wire \EXU/_1138_ ;
wire \EXU/_1139_ ;
wire \EXU/_1140_ ;
wire \EXU/_1141_ ;
wire \EXU/_1142_ ;
wire \EXU/_1143_ ;
wire \EXU/_1144_ ;
wire \EXU/_1145_ ;
wire \EXU/_1146_ ;
wire \EXU/_1147_ ;
wire \EXU/_1148_ ;
wire \EXU/_1149_ ;
wire \EXU/_1150_ ;
wire \EXU/_1151_ ;
wire \EXU/_1152_ ;
wire \EXU/_1153_ ;
wire \EXU/_1154_ ;
wire \EXU/_1155_ ;
wire \EXU/_1156_ ;
wire \EXU/_1157_ ;
wire \EXU/_1158_ ;
wire \EXU/_1159_ ;
wire \EXU/_1160_ ;
wire \EXU/_1161_ ;
wire \EXU/_1162_ ;
wire \EXU/_1163_ ;
wire \EXU/_1164_ ;
wire \EXU/_1165_ ;
wire \EXU/_1166_ ;
wire \EXU/_1167_ ;
wire \EXU/_1168_ ;
wire \EXU/_1169_ ;
wire \EXU/_1170_ ;
wire \EXU/_1171_ ;
wire \EXU/_1172_ ;
wire \EXU/_1173_ ;
wire \EXU/_1174_ ;
wire \EXU/_1175_ ;
wire \EXU/_1176_ ;
wire \EXU/_1177_ ;
wire \EXU/_1178_ ;
wire \EXU/_1179_ ;
wire \EXU/_1180_ ;
wire \EXU/_1181_ ;
wire \EXU/_1182_ ;
wire \EXU/_1183_ ;
wire \EXU/_1184_ ;
wire \EXU/_1185_ ;
wire \EXU/_1186_ ;
wire \EXU/_1187_ ;
wire \EXU/_1188_ ;
wire \EXU/_1189_ ;
wire \EXU/_1190_ ;
wire \EXU/_1191_ ;
wire \EXU/_1192_ ;
wire \EXU/_1193_ ;
wire \EXU/_1194_ ;
wire \EXU/_1195_ ;
wire \EXU/_1196_ ;
wire \EXU/_1197_ ;
wire \EXU/_1198_ ;
wire \EXU/_1199_ ;
wire \EXU/_1200_ ;
wire \EXU/_1201_ ;
wire \EXU/_1202_ ;
wire \EXU/_1203_ ;
wire \EXU/_1204_ ;
wire \EXU/_1205_ ;
wire \EXU/_1206_ ;
wire \EXU/_1207_ ;
wire \EXU/_1208_ ;
wire \EXU/_1209_ ;
wire \EXU/_1210_ ;
wire \EXU/_1211_ ;
wire \EXU/_1212_ ;
wire \EXU/_1213_ ;
wire \EXU/_1214_ ;
wire \EXU/_1215_ ;
wire \EXU/_1216_ ;
wire \EXU/_1217_ ;
wire \EXU/_1218_ ;
wire \EXU/_1219_ ;
wire \EXU/_1220_ ;
wire \EXU/_1221_ ;
wire \EXU/_1222_ ;
wire \EXU/_1223_ ;
wire \EXU/_1224_ ;
wire \EXU/_1225_ ;
wire \EXU/_1226_ ;
wire \EXU/_1227_ ;
wire \EXU/_1228_ ;
wire \EXU/_1229_ ;
wire \EXU/_1230_ ;
wire \EXU/_1231_ ;
wire \EXU/_1232_ ;
wire \EXU/_1233_ ;
wire \EXU/_1234_ ;
wire \EXU/_1235_ ;
wire \EXU/_1236_ ;
wire \EXU/_1237_ ;
wire \EXU/_1238_ ;
wire \EXU/_1239_ ;
wire \EXU/_1240_ ;
wire \EXU/_1241_ ;
wire \EXU/_1242_ ;
wire \EXU/_1243_ ;
wire \EXU/_1244_ ;
wire \EXU/_1245_ ;
wire \EXU/_1246_ ;
wire \EXU/_1247_ ;
wire \EXU/_1248_ ;
wire \EXU/_1249_ ;
wire \EXU/_1250_ ;
wire \EXU/_1251_ ;
wire \EXU/_1252_ ;
wire \EXU/_1253_ ;
wire \EXU/_1254_ ;
wire \EXU/_1255_ ;
wire \EXU/_1256_ ;
wire \EXU/_1257_ ;
wire \EXU/_1258_ ;
wire \EXU/_1259_ ;
wire \EXU/_1260_ ;
wire \EXU/_1261_ ;
wire \EXU/_1262_ ;
wire \EXU/_1263_ ;
wire \EXU/_1264_ ;
wire \EXU/_1265_ ;
wire \EXU/_1266_ ;
wire \EXU/_1267_ ;
wire \EXU/_1268_ ;
wire \EXU/_1269_ ;
wire \EXU/_1270_ ;
wire \EXU/_1271_ ;
wire \EXU/_1272_ ;
wire \EXU/_1273_ ;
wire \EXU/_1274_ ;
wire \EXU/_1275_ ;
wire \EXU/_1276_ ;
wire \EXU/_1277_ ;
wire \EXU/_1278_ ;
wire \EXU/_1279_ ;
wire \EXU/_1280_ ;
wire \EXU/_1281_ ;
wire \EXU/_1282_ ;
wire \EXU/_1283_ ;
wire \EXU/_1284_ ;
wire \EXU/_1285_ ;
wire \EXU/_1286_ ;
wire \EXU/_1287_ ;
wire \EXU/_1288_ ;
wire \EXU/_1289_ ;
wire \EXU/_1290_ ;
wire \EXU/_1291_ ;
wire \EXU/_1292_ ;
wire \EXU/_1293_ ;
wire \EXU/_1294_ ;
wire \EXU/_1295_ ;
wire \EXU/_1296_ ;
wire \EXU/_1297_ ;
wire \EXU/_1298_ ;
wire \EXU/_1299_ ;
wire \EXU/_1300_ ;
wire \EXU/_1301_ ;
wire \EXU/_1302_ ;
wire \EXU/_1303_ ;
wire \EXU/_1304_ ;
wire \EXU/_1305_ ;
wire \EXU/_1306_ ;
wire \EXU/_1307_ ;
wire \EXU/_1308_ ;
wire \EXU/_1309_ ;
wire \EXU/_1310_ ;
wire \EXU/_1311_ ;
wire \EXU/_1312_ ;
wire \EXU/_1313_ ;
wire \EXU/_1314_ ;
wire \EXU/_1315_ ;
wire \EXU/_1316_ ;
wire \EXU/_1317_ ;
wire \EXU/_1318_ ;
wire \EXU/_1319_ ;
wire \EXU/_1320_ ;
wire \EXU/_1321_ ;
wire \EXU/_1322_ ;
wire \EXU/_1323_ ;
wire \EXU/_1324_ ;
wire \EXU/_1325_ ;
wire \EXU/_1326_ ;
wire \EXU/_1327_ ;
wire \EXU/_1328_ ;
wire \EXU/_1329_ ;
wire \EXU/_1330_ ;
wire \EXU/_1331_ ;
wire \EXU/_1332_ ;
wire \EXU/_1333_ ;
wire \EXU/_1334_ ;
wire \EXU/_1335_ ;
wire \EXU/_1336_ ;
wire \EXU/_1337_ ;
wire \EXU/_1338_ ;
wire \EXU/_1339_ ;
wire \EXU/_1340_ ;
wire \EXU/_1341_ ;
wire \EXU/_1342_ ;
wire \EXU/_1343_ ;
wire \EXU/_1344_ ;
wire \EXU/_1345_ ;
wire \EXU/_1346_ ;
wire \EXU/_1347_ ;
wire \EXU/_1348_ ;
wire \EXU/_1349_ ;
wire \EXU/_1350_ ;
wire \EXU/_1351_ ;
wire \EXU/_1352_ ;
wire \EXU/_1353_ ;
wire \EXU/_1354_ ;
wire \EXU/_1355_ ;
wire \EXU/_1356_ ;
wire \EXU/_1357_ ;
wire \EXU/_1358_ ;
wire \EXU/_1359_ ;
wire \EXU/_1360_ ;
wire \EXU/_1361_ ;
wire \EXU/_1362_ ;
wire \EXU/_1363_ ;
wire \EXU/_1364_ ;
wire \EXU/_1365_ ;
wire \EXU/_1366_ ;
wire \EXU/_1367_ ;
wire \EXU/_1368_ ;
wire \EXU/_1369_ ;
wire \EXU/_1370_ ;
wire \EXU/_1371_ ;
wire \EXU/_1372_ ;
wire \EXU/_1373_ ;
wire \EXU/_1374_ ;
wire \EXU/_1375_ ;
wire \EXU/_1376_ ;
wire \EXU/_1377_ ;
wire \EXU/_1378_ ;
wire \EXU/_1379_ ;
wire \EXU/_1380_ ;
wire \EXU/_1381_ ;
wire \EXU/_1382_ ;
wire \EXU/_1383_ ;
wire \EXU/_1384_ ;
wire \EXU/_1385_ ;
wire \EXU/_1386_ ;
wire \EXU/_1387_ ;
wire \EXU/_1388_ ;
wire \EXU/_1389_ ;
wire \EXU/_1390_ ;
wire \EXU/_1391_ ;
wire \EXU/_1392_ ;
wire \EXU/_1393_ ;
wire \EXU/_1394_ ;
wire \EXU/_1395_ ;
wire \EXU/_1396_ ;
wire \EXU/_1397_ ;
wire \EXU/_1398_ ;
wire \EXU/_1399_ ;
wire \EXU/_1400_ ;
wire \EXU/_1401_ ;
wire \EXU/_1402_ ;
wire \EXU/_1403_ ;
wire \EXU/_1404_ ;
wire \EXU/_1405_ ;
wire \EXU/_1406_ ;
wire \EXU/_1407_ ;
wire \EXU/_1408_ ;
wire \EXU/_1409_ ;
wire \EXU/_1410_ ;
wire \EXU/_1411_ ;
wire \EXU/_1412_ ;
wire \EXU/_1413_ ;
wire \EXU/_1414_ ;
wire \EXU/_1415_ ;
wire \EXU/_1416_ ;
wire \EXU/_1417_ ;
wire \EXU/_1418_ ;
wire \EXU/_1419_ ;
wire \EXU/_1420_ ;
wire \EXU/_1421_ ;
wire \EXU/_1422_ ;
wire \EXU/_1423_ ;
wire \EXU/_1424_ ;
wire \EXU/_1425_ ;
wire \EXU/_1426_ ;
wire \EXU/_1427_ ;
wire \EXU/_1428_ ;
wire \EXU/_1429_ ;
wire \EXU/_1430_ ;
wire \EXU/_1431_ ;
wire \EXU/_1432_ ;
wire \EXU/_1433_ ;
wire \EXU/_1434_ ;
wire \EXU/_1435_ ;
wire \EXU/_1436_ ;
wire \EXU/_1437_ ;
wire \EXU/_1438_ ;
wire \EXU/_1439_ ;
wire \EXU/_1440_ ;
wire \EXU/_1441_ ;
wire \EXU/_1442_ ;
wire \EXU/_1443_ ;
wire \EXU/_1444_ ;
wire \EXU/_1445_ ;
wire \EXU/_1446_ ;
wire \EXU/_1447_ ;
wire \EXU/_1448_ ;
wire \EXU/_1449_ ;
wire \EXU/_1450_ ;
wire \EXU/_1451_ ;
wire \EXU/_1452_ ;
wire \EXU/_1453_ ;
wire \EXU/_1454_ ;
wire \EXU/_1455_ ;
wire \EXU/_1456_ ;
wire \EXU/_1457_ ;
wire \EXU/_1458_ ;
wire \EXU/_1459_ ;
wire \EXU/_1460_ ;
wire \EXU/_1461_ ;
wire \EXU/_1462_ ;
wire \EXU/_1463_ ;
wire \EXU/_1464_ ;
wire \EXU/_1465_ ;
wire \EXU/_1466_ ;
wire \EXU/_1467_ ;
wire \EXU/_1468_ ;
wire \EXU/_1469_ ;
wire \EXU/_1470_ ;
wire \EXU/_1471_ ;
wire \EXU/_1472_ ;
wire \EXU/_1473_ ;
wire \EXU/_1474_ ;
wire \EXU/_1475_ ;
wire \EXU/_1476_ ;
wire \EXU/_1477_ ;
wire \EXU/_1478_ ;
wire \EXU/_1479_ ;
wire \EXU/_1480_ ;
wire \EXU/_1481_ ;
wire \EXU/_1482_ ;
wire \EXU/_1483_ ;
wire \EXU/_1484_ ;
wire \EXU/_1485_ ;
wire \EXU/_1486_ ;
wire \EXU/_1487_ ;
wire \EXU/_1488_ ;
wire \EXU/_1489_ ;
wire \EXU/_1490_ ;
wire \EXU/_1491_ ;
wire \EXU/_1492_ ;
wire \EXU/_1493_ ;
wire \EXU/_1494_ ;
wire \EXU/_1495_ ;
wire \EXU/_1496_ ;
wire \EXU/_1497_ ;
wire \EXU/_1498_ ;
wire \EXU/_1499_ ;
wire \EXU/_1500_ ;
wire \EXU/_1501_ ;
wire \EXU/_1502_ ;
wire \EXU/_1503_ ;
wire \EXU/_1504_ ;
wire \EXU/_1505_ ;
wire \EXU/_1506_ ;
wire \EXU/_1507_ ;
wire \EXU/_1508_ ;
wire \EXU/_1509_ ;
wire \EXU/_1510_ ;
wire \EXU/_1511_ ;
wire \EXU/_1512_ ;
wire \EXU/_1513_ ;
wire \EXU/_1514_ ;
wire \EXU/_1515_ ;
wire \EXU/_1516_ ;
wire \EXU/_1517_ ;
wire \EXU/_1518_ ;
wire \EXU/_1519_ ;
wire \EXU/_1520_ ;
wire \EXU/_1521_ ;
wire \EXU/_1522_ ;
wire \EXU/_1523_ ;
wire \EXU/_1524_ ;
wire \EXU/_1525_ ;
wire \EXU/_1526_ ;
wire \EXU/_1527_ ;
wire \EXU/_1528_ ;
wire \EXU/_1529_ ;
wire \EXU/_1530_ ;
wire \EXU/_1531_ ;
wire \EXU/_1532_ ;
wire \EXU/_1533_ ;
wire \EXU/_1534_ ;
wire \EXU/_1535_ ;
wire \EXU/_1536_ ;
wire \EXU/_1537_ ;
wire \EXU/_1538_ ;
wire \EXU/_1539_ ;
wire \EXU/_1540_ ;
wire \EXU/_1541_ ;
wire \EXU/_1542_ ;
wire \EXU/_1543_ ;
wire \EXU/_1544_ ;
wire \EXU/_1545_ ;
wire \EXU/_1546_ ;
wire \EXU/_1547_ ;
wire \EXU/_1548_ ;
wire \EXU/_1549_ ;
wire \EXU/_1550_ ;
wire \EXU/_1551_ ;
wire \EXU/_1552_ ;
wire \EXU/_1553_ ;
wire \EXU/_1554_ ;
wire \EXU/_1555_ ;
wire \EXU/_1556_ ;
wire \EXU/_1557_ ;
wire \EXU/_1558_ ;
wire \EXU/_1559_ ;
wire \EXU/_1560_ ;
wire \EXU/_1561_ ;
wire \EXU/_1562_ ;
wire \EXU/_1563_ ;
wire \EXU/_1564_ ;
wire \EXU/_1565_ ;
wire \EXU/_1566_ ;
wire \EXU/_1567_ ;
wire \EXU/_1568_ ;
wire \EXU/_1569_ ;
wire \EXU/_1570_ ;
wire \EXU/_1571_ ;
wire \EXU/_1572_ ;
wire \EXU/_1573_ ;
wire \EXU/_1574_ ;
wire \EXU/_1575_ ;
wire \EXU/_1576_ ;
wire \EXU/_1577_ ;
wire \EXU/_1578_ ;
wire \EXU/_1579_ ;
wire \EXU/_1580_ ;
wire \EXU/_1581_ ;
wire \EXU/_1582_ ;
wire \EXU/_1583_ ;
wire \EXU/_1584_ ;
wire \EXU/_1585_ ;
wire \EXU/_1586_ ;
wire \EXU/_1587_ ;
wire \EXU/_1588_ ;
wire \EXU/_1589_ ;
wire \EXU/_1590_ ;
wire \EXU/_1591_ ;
wire \EXU/_1592_ ;
wire \EXU/_1593_ ;
wire \EXU/_1594_ ;
wire \EXU/_1595_ ;
wire \EXU/_1596_ ;
wire \EXU/_1597_ ;
wire \EXU/_1598_ ;
wire \EXU/_1599_ ;
wire \EXU/_1600_ ;
wire \EXU/_1601_ ;
wire \EXU/_1602_ ;
wire \EXU/_1603_ ;
wire \EXU/_1604_ ;
wire \EXU/_1605_ ;
wire \EXU/_1606_ ;
wire \EXU/_1607_ ;
wire \EXU/_1608_ ;
wire \EXU/_1609_ ;
wire \EXU/_1610_ ;
wire \EXU/_1611_ ;
wire \EXU/_1612_ ;
wire \EXU/_1613_ ;
wire \EXU/_1614_ ;
wire \EXU/_1615_ ;
wire \EXU/_1616_ ;
wire \EXU/_1617_ ;
wire \EXU/_1618_ ;
wire \EXU/_1619_ ;
wire \EXU/_1620_ ;
wire \EXU/_1621_ ;
wire \EXU/_1622_ ;
wire \EXU/_1623_ ;
wire \EXU/_1624_ ;
wire \EXU/_1625_ ;
wire \EXU/_1626_ ;
wire \EXU/_1627_ ;
wire \EXU/_1628_ ;
wire \EXU/_1629_ ;
wire \EXU/_1630_ ;
wire \EXU/_1631_ ;
wire \EXU/_1632_ ;
wire \EXU/_1633_ ;
wire \EXU/_1634_ ;
wire \EXU/_1635_ ;
wire \EXU/_1636_ ;
wire \EXU/_1637_ ;
wire \EXU/_1638_ ;
wire \EXU/_1639_ ;
wire \EXU/_1640_ ;
wire \EXU/_1641_ ;
wire \EXU/_1642_ ;
wire \EXU/_ALU_io_less ;
wire \EXU/_ALU_io_zero ;
wire \EXU/_BrCond_io_PCASrc ;
wire \EXU/_BrCond_io_PCBSrc ;
wire \EXU/in_control_aluASrc ;
wire \EXU/in_control_csrSrc ;
wire \EXU/ALU/_000_ ;
wire \EXU/ALU/_001_ ;
wire \EXU/ALU/_002_ ;
wire \EXU/ALU/_003_ ;
wire \EXU/ALU/_004_ ;
wire \EXU/ALU/_005_ ;
wire \EXU/ALU/_006_ ;
wire \EXU/ALU/_007_ ;
wire \EXU/ALU/_008_ ;
wire \EXU/ALU/_009_ ;
wire \EXU/ALU/_010_ ;
wire \EXU/ALU/_011_ ;
wire \EXU/ALU/_012_ ;
wire \EXU/ALU/_013_ ;
wire \EXU/ALU/_014_ ;
wire \EXU/ALU/_015_ ;
wire \EXU/ALU/_016_ ;
wire \EXU/ALU/_017_ ;
wire \EXU/ALU/_018_ ;
wire \EXU/ALU/_019_ ;
wire \EXU/ALU/_020_ ;
wire \EXU/ALU/_021_ ;
wire \EXU/ALU/_022_ ;
wire \EXU/ALU/_023_ ;
wire \EXU/ALU/_024_ ;
wire \EXU/ALU/_025_ ;
wire \EXU/ALU/_026_ ;
wire \EXU/ALU/_027_ ;
wire \EXU/ALU/_028_ ;
wire \EXU/ALU/_029_ ;
wire \EXU/ALU/_030_ ;
wire \EXU/ALU/_031_ ;
wire \EXU/ALU/_032_ ;
wire \EXU/ALU/_033_ ;
wire \EXU/ALU/_034_ ;
wire \EXU/ALU/_035_ ;
wire \EXU/ALU/_036_ ;
wire \EXU/ALU/_037_ ;
wire \EXU/ALU/_038_ ;
wire \EXU/ALU/_039_ ;
wire \EXU/ALU/_040_ ;
wire \EXU/ALU/_041_ ;
wire \EXU/ALU/_042_ ;
wire \EXU/ALU/_043_ ;
wire \EXU/ALU/_044_ ;
wire \EXU/ALU/_045_ ;
wire \EXU/ALU/_046_ ;
wire \EXU/ALU/_047_ ;
wire \EXU/ALU/_048_ ;
wire \EXU/ALU/_049_ ;
wire \EXU/ALU/_050_ ;
wire \EXU/ALU/_051_ ;
wire \EXU/ALU/_052_ ;
wire \EXU/ALU/_053_ ;
wire \EXU/ALU/_054_ ;
wire \EXU/ALU/_055_ ;
wire \EXU/ALU/_056_ ;
wire \EXU/ALU/_057_ ;
wire \EXU/ALU/_058_ ;
wire \EXU/ALU/_059_ ;
wire \EXU/ALU/_060_ ;
wire \EXU/ALU/_061_ ;
wire \EXU/ALU/_062_ ;
wire \EXU/ALU/_063_ ;
wire \EXU/ALU/_064_ ;
wire \EXU/ALU/_065_ ;
wire \EXU/ALU/_066_ ;
wire \EXU/ALU/_067_ ;
wire \EXU/ALU/_068_ ;
wire \EXU/ALU/_069_ ;
wire \EXU/ALU/_070_ ;
wire \EXU/ALU/_071_ ;
wire \EXU/ALU/_072_ ;
wire \EXU/ALU/_073_ ;
wire \EXU/ALU/_074_ ;
wire \EXU/ALU/_075_ ;
wire \EXU/ALU/_076_ ;
wire \EXU/ALU/_077_ ;
wire \EXU/ALU/_078_ ;
wire \EXU/ALU/_079_ ;
wire \EXU/ALU/_080_ ;
wire \EXU/ALU/_081_ ;
wire \EXU/ALU/_082_ ;
wire \EXU/ALU/_083_ ;
wire \EXU/ALU/_084_ ;
wire \EXU/ALU/_085_ ;
wire \EXU/ALU/_086_ ;
wire \EXU/ALU/_087_ ;
wire \EXU/ALU/_088_ ;
wire \EXU/ALU/_089_ ;
wire \EXU/ALU/_090_ ;
wire \EXU/ALU/_091_ ;
wire \EXU/ALU/_092_ ;
wire \EXU/ALU/_093_ ;
wire \EXU/ALU/_094_ ;
wire \EXU/ALU/_095_ ;
wire \EXU/ALU/_096_ ;
wire \EXU/ALU/_097_ ;
wire \EXU/ALU/_098_ ;
wire \EXU/ALU/_099_ ;
wire \EXU/ALU/_100_ ;
wire \EXU/ALU/_101_ ;
wire \EXU/ALU/_102_ ;
wire \EXU/ALU/_103_ ;
wire \EXU/ALU/_104_ ;
wire \EXU/ALU/_105_ ;
wire \EXU/ALU/_106_ ;
wire \EXU/ALU/_107_ ;
wire \EXU/ALU/_108_ ;
wire \EXU/ALU/_109_ ;
wire \EXU/ALU/_110_ ;
wire \EXU/ALU/_111_ ;
wire \EXU/ALU/_112_ ;
wire \EXU/ALU/_113_ ;
wire \EXU/ALU/_114_ ;
wire \EXU/ALU/_115_ ;
wire \EXU/ALU/_116_ ;
wire \EXU/ALU/_117_ ;
wire \EXU/ALU/_118_ ;
wire \EXU/ALU/_119_ ;
wire \EXU/ALU/_120_ ;
wire \EXU/ALU/_121_ ;
wire \EXU/ALU/_122_ ;
wire \EXU/ALU/_123_ ;
wire \EXU/ALU/_124_ ;
wire \EXU/ALU/_125_ ;
wire \EXU/ALU/_126_ ;
wire \EXU/ALU/_127_ ;
wire \EXU/ALU/_128_ ;
wire \EXU/ALU/_129_ ;
wire \EXU/ALU/_130_ ;
wire \EXU/ALU/_131_ ;
wire \EXU/ALU/_132_ ;
wire \EXU/ALU/_133_ ;
wire \EXU/ALU/_134_ ;
wire \EXU/ALU/_135_ ;
wire \EXU/ALU/_136_ ;
wire \EXU/ALU/_137_ ;
wire \EXU/ALU/_138_ ;
wire \EXU/ALU/_139_ ;
wire \EXU/ALU/_140_ ;
wire \EXU/ALU/_141_ ;
wire \EXU/ALU/_142_ ;
wire \EXU/ALU/_143_ ;
wire \EXU/ALU/_144_ ;
wire \EXU/ALU/_145_ ;
wire \EXU/ALU/_146_ ;
wire \EXU/ALU/_147_ ;
wire \EXU/ALU/_148_ ;
wire \EXU/ALU/_149_ ;
wire \EXU/ALU/_150_ ;
wire \EXU/ALU/_151_ ;
wire \EXU/ALU/_152_ ;
wire \EXU/ALU/_153_ ;
wire \EXU/ALU/_154_ ;
wire \EXU/ALU/_155_ ;
wire \EXU/ALU/_156_ ;
wire \EXU/ALU/_157_ ;
wire \EXU/ALU/_158_ ;
wire \EXU/ALU/_159_ ;
wire \EXU/ALU/_160_ ;
wire \EXU/ALU/_161_ ;
wire \EXU/ALU/_162_ ;
wire \EXU/ALU/_163_ ;
wire \EXU/ALU/_164_ ;
wire \EXU/ALU/_165_ ;
wire \EXU/ALU/_166_ ;
wire \EXU/ALU/_167_ ;
wire \EXU/ALU/_168_ ;
wire \EXU/ALU/_169_ ;
wire \EXU/ALU/_170_ ;
wire \EXU/ALU/_171_ ;
wire \EXU/ALU/_172_ ;
wire \EXU/ALU/_173_ ;
wire \EXU/ALU/_174_ ;
wire \EXU/ALU/_175_ ;
wire \EXU/ALU/_176_ ;
wire \EXU/ALU/_177_ ;
wire \EXU/ALU/_178_ ;
wire \EXU/ALU/_179_ ;
wire \EXU/ALU/_180_ ;
wire \EXU/ALU/_181_ ;
wire \EXU/ALU/_182_ ;
wire \EXU/ALU/_183_ ;
wire \EXU/ALU/_184_ ;
wire \EXU/ALU/_185_ ;
wire \EXU/ALU/_186_ ;
wire \EXU/ALU/_187_ ;
wire \EXU/ALU/_188_ ;
wire \EXU/ALU/_189_ ;
wire \EXU/ALU/_190_ ;
wire \EXU/ALU/_191_ ;
wire \EXU/ALU/_192_ ;
wire \EXU/ALU/_193_ ;
wire \EXU/ALU/_194_ ;
wire \EXU/ALU/_195_ ;
wire \EXU/ALU/_196_ ;
wire \EXU/ALU/_197_ ;
wire \EXU/ALU/_198_ ;
wire \EXU/ALU/_199_ ;
wire \EXU/ALU/_200_ ;
wire \EXU/ALU/_201_ ;
wire \EXU/ALU/_202_ ;
wire \EXU/ALU/_203_ ;
wire \EXU/ALU/_204_ ;
wire \EXU/ALU/_205_ ;
wire \EXU/ALU/_206_ ;
wire \EXU/ALU/_207_ ;
wire \EXU/ALU/_208_ ;
wire \EXU/ALU/_209_ ;
wire \EXU/ALU/_210_ ;
wire \EXU/ALU/_211_ ;
wire \EXU/ALU/_212_ ;
wire \EXU/ALU/_213_ ;
wire \EXU/ALU/_214_ ;
wire \EXU/ALU/_215_ ;
wire \EXU/ALU/_216_ ;
wire \EXU/ALU/_217_ ;
wire \EXU/ALU/_218_ ;
wire \EXU/ALU/_219_ ;
wire \EXU/ALU/_220_ ;
wire \EXU/ALU/_221_ ;
wire \EXU/ALU/_222_ ;
wire \EXU/ALU/_223_ ;
wire \EXU/ALU/_224_ ;
wire \EXU/ALU/_225_ ;
wire \EXU/ALU/_226_ ;
wire \EXU/ALU/_227_ ;
wire \EXU/ALU/_228_ ;
wire \EXU/ALU/_229_ ;
wire \EXU/ALU/_230_ ;
wire \EXU/ALU/_231_ ;
wire \EXU/ALU/_232_ ;
wire \EXU/ALU/_233_ ;
wire \EXU/ALU/_234_ ;
wire \EXU/ALU/_235_ ;
wire \EXU/ALU/_236_ ;
wire \EXU/ALU/_237_ ;
wire \EXU/ALU/_238_ ;
wire \EXU/ALU/_239_ ;
wire \EXU/ALU/_240_ ;
wire \EXU/ALU/_241_ ;
wire \EXU/ALU/_242_ ;
wire \EXU/ALU/_243_ ;
wire \EXU/ALU/_244_ ;
wire \EXU/ALU/_245_ ;
wire \EXU/ALU/_246_ ;
wire \EXU/ALU/_247_ ;
wire \EXU/ALU/_248_ ;
wire \EXU/ALU/_249_ ;
wire \EXU/ALU/_250_ ;
wire \EXU/ALU/_251_ ;
wire \EXU/ALU/_252_ ;
wire \EXU/ALU/_253_ ;
wire \EXU/ALU/_254_ ;
wire \EXU/ALU/_255_ ;
wire \EXU/ALU/_256_ ;
wire \EXU/ALU/_257_ ;
wire \EXU/ALU/_258_ ;
wire \EXU/ALU/_259_ ;
wire \EXU/ALU/_260_ ;
wire \EXU/ALU/_261_ ;
wire \EXU/ALU/_262_ ;
wire \EXU/ALU/_263_ ;
wire \EXU/ALU/_264_ ;
wire \EXU/ALU/_265_ ;
wire \EXU/ALU/_266_ ;
wire \EXU/ALU/_267_ ;
wire \EXU/ALU/_268_ ;
wire \EXU/ALU/_269_ ;
wire \EXU/ALU/_270_ ;
wire \EXU/ALU/_271_ ;
wire \EXU/ALU/_272_ ;
wire \EXU/ALU/_273_ ;
wire \EXU/ALU/_274_ ;
wire \EXU/ALU/_275_ ;
wire \EXU/ALU/_276_ ;
wire \EXU/ALU/_277_ ;
wire \EXU/ALU/_278_ ;
wire \EXU/ALU/_279_ ;
wire \EXU/ALU/_280_ ;
wire \EXU/ALU/_281_ ;
wire \EXU/ALU/_282_ ;
wire \EXU/ALU/_283_ ;
wire \EXU/ALU/_284_ ;
wire \EXU/ALU/_285_ ;
wire \EXU/ALU/_286_ ;
wire \EXU/ALU/_287_ ;
wire \EXU/ALU/_288_ ;
wire \EXU/ALU/_289_ ;
wire \EXU/ALU/_290_ ;
wire \EXU/ALU/_291_ ;
wire \EXU/ALU/_292_ ;
wire \EXU/ALU/_293_ ;
wire \EXU/ALU/_294_ ;
wire \EXU/ALU/_295_ ;
wire \EXU/ALU/_296_ ;
wire \EXU/ALU/_297_ ;
wire \EXU/ALU/_298_ ;
wire \EXU/ALU/_299_ ;
wire \EXU/ALU/_300_ ;
wire \EXU/ALU/_301_ ;
wire \EXU/ALU/_302_ ;
wire \EXU/ALU/_303_ ;
wire \EXU/ALU/_304_ ;
wire \EXU/ALU/_305_ ;
wire \EXU/ALU/_306_ ;
wire \EXU/ALU/_307_ ;
wire \EXU/ALU/_308_ ;
wire \EXU/ALU/_309_ ;
wire \EXU/ALU/_310_ ;
wire \EXU/ALU/_311_ ;
wire \EXU/ALU/_312_ ;
wire \EXU/ALU/_313_ ;
wire \EXU/ALU/_314_ ;
wire \EXU/ALU/_315_ ;
wire \EXU/ALU/_316_ ;
wire \EXU/ALU/_317_ ;
wire \EXU/ALU/_318_ ;
wire \EXU/ALU/_319_ ;
wire \EXU/ALU/_320_ ;
wire \EXU/ALU/_321_ ;
wire \EXU/ALU/_322_ ;
wire \EXU/ALU/_323_ ;
wire \EXU/ALU/_324_ ;
wire \EXU/ALU/_325_ ;
wire \EXU/ALU/_326_ ;
wire \EXU/ALU/_327_ ;
wire \EXU/ALU/_328_ ;
wire \EXU/ALU/_329_ ;
wire \EXU/ALU/_330_ ;
wire \EXU/ALU/_331_ ;
wire \EXU/ALU/_332_ ;
wire \EXU/ALU/_333_ ;
wire \EXU/ALU/_334_ ;
wire \EXU/ALU/_335_ ;
wire \EXU/ALU/_336_ ;
wire \EXU/ALU/_337_ ;
wire \EXU/ALU/_338_ ;
wire \EXU/ALU/_339_ ;
wire \EXU/ALU/_340_ ;
wire \EXU/ALU/_341_ ;
wire \EXU/ALU/_342_ ;
wire \EXU/ALU/_343_ ;
wire \EXU/ALU/_344_ ;
wire \EXU/ALU/_345_ ;
wire \EXU/ALU/_346_ ;
wire \EXU/ALU/_347_ ;
wire \EXU/ALU/_348_ ;
wire \EXU/ALU/_349_ ;
wire \EXU/ALU/_350_ ;
wire \EXU/ALU/_351_ ;
wire \EXU/ALU/_352_ ;
wire \EXU/ALU/_353_ ;
wire \EXU/ALU/_354_ ;
wire \EXU/ALU/_355_ ;
wire \EXU/ALU/_356_ ;
wire \EXU/ALU/_357_ ;
wire \EXU/ALU/_358_ ;
wire \EXU/ALU/_359_ ;
wire \EXU/ALU/_360_ ;
wire \EXU/ALU/_361_ ;
wire \EXU/ALU/_362_ ;
wire \EXU/ALU/_363_ ;
wire \EXU/ALU/_364_ ;
wire \EXU/ALU/_365_ ;
wire \EXU/ALU/_366_ ;
wire \EXU/ALU/_367_ ;
wire \EXU/ALU/_368_ ;
wire \EXU/ALU/_369_ ;
wire \EXU/ALU/_370_ ;
wire \EXU/ALU/_371_ ;
wire \EXU/ALU/_372_ ;
wire \EXU/ALU/_373_ ;
wire \EXU/ALU/_374_ ;
wire \EXU/ALU/_375_ ;
wire \EXU/ALU/_376_ ;
wire \EXU/ALU/_377_ ;
wire \EXU/ALU/_378_ ;
wire \EXU/ALU/_379_ ;
wire \EXU/ALU/_380_ ;
wire \EXU/ALU/_381_ ;
wire \EXU/ALU/_382_ ;
wire \EXU/ALU/_383_ ;
wire \EXU/ALU/_384_ ;
wire \EXU/ALU/_385_ ;
wire \EXU/ALU/_386_ ;
wire \EXU/ALU/_387_ ;
wire \EXU/ALU/_388_ ;
wire \EXU/ALU/_389_ ;
wire \EXU/ALU/_390_ ;
wire \EXU/ALU/_391_ ;
wire \EXU/ALU/_392_ ;
wire \EXU/ALU/_393_ ;
wire \EXU/ALU/_394_ ;
wire \EXU/ALU/_395_ ;
wire \EXU/ALU/_396_ ;
wire \EXU/ALU/_397_ ;
wire \EXU/ALU/_398_ ;
wire \EXU/ALU/_399_ ;
wire \EXU/ALU/_400_ ;
wire \EXU/ALU/_401_ ;
wire \EXU/ALU/_402_ ;
wire \EXU/ALU/_403_ ;
wire \EXU/ALU/_404_ ;
wire \EXU/ALU/_405_ ;
wire \EXU/ALU/_406_ ;
wire \EXU/ALU/_407_ ;
wire \EXU/ALU/_408_ ;
wire \EXU/ALU/_409_ ;
wire \EXU/ALU/_410_ ;
wire \EXU/ALU/_411_ ;
wire \EXU/ALU/_412_ ;
wire \EXU/ALU/_413_ ;
wire \EXU/ALU/_414_ ;
wire \EXU/ALU/_415_ ;
wire \EXU/ALU/_416_ ;
wire \EXU/ALU/_417_ ;
wire \EXU/ALU/_418_ ;
wire \EXU/ALU/_419_ ;
wire \EXU/ALU/_420_ ;
wire \EXU/ALU/_421_ ;
wire \EXU/ALU/_422_ ;
wire \EXU/ALU/_423_ ;
wire \EXU/ALU/_424_ ;
wire \EXU/ALU/_425_ ;
wire \EXU/ALU/_426_ ;
wire \EXU/ALU/_427_ ;
wire \EXU/ALU/_428_ ;
wire \EXU/ALU/_429_ ;
wire \EXU/ALU/_430_ ;
wire \EXU/ALU/_431_ ;
wire \EXU/ALU/_432_ ;
wire \EXU/ALU/_433_ ;
wire \EXU/ALU/_434_ ;
wire \EXU/ALU/_435_ ;
wire \EXU/ALU/_436_ ;
wire \EXU/ALU/_437_ ;
wire \EXU/ALU/_438_ ;
wire \EXU/ALU/_439_ ;
wire \EXU/ALU/_440_ ;
wire \EXU/ALU/_441_ ;
wire \EXU/ALU/_442_ ;
wire \EXU/ALU/_443_ ;
wire \EXU/ALU/_444_ ;
wire \EXU/ALU/_445_ ;
wire \EXU/ALU/_446_ ;
wire \EXU/ALU/_447_ ;
wire \EXU/ALU/_448_ ;
wire \EXU/ALU/_449_ ;
wire \EXU/ALU/_450_ ;
wire \EXU/ALU/_451_ ;
wire \EXU/ALU/_452_ ;
wire \EXU/ALU/_453_ ;
wire \EXU/ALU/_454_ ;
wire \EXU/ALU/_455_ ;
wire \EXU/ALU/_456_ ;
wire \EXU/ALU/_457_ ;
wire \EXU/ALU/_adder_io_carry ;
wire \EXU/ALU/_adder_io_overflow ;
wire \EXU/ALU/_aluControl_io_isArith ;
wire \EXU/ALU/_aluControl_io_isLeft ;
wire \EXU/ALU/_aluControl_io_isSub ;
wire \EXU/ALU/_aluControl_io_isUnsigned ;
wire \EXU/ALU/adder/_000_ ;
wire \EXU/ALU/adder/_001_ ;
wire \EXU/ALU/adder/_002_ ;
wire \EXU/ALU/adder/_003_ ;
wire \EXU/ALU/adder/_004_ ;
wire \EXU/ALU/adder/_005_ ;
wire \EXU/ALU/adder/_006_ ;
wire \EXU/ALU/adder/_007_ ;
wire \EXU/ALU/adder/_008_ ;
wire \EXU/ALU/adder/_009_ ;
wire \EXU/ALU/adder/_010_ ;
wire \EXU/ALU/adder/_011_ ;
wire \EXU/ALU/adder/_012_ ;
wire \EXU/ALU/adder/_013_ ;
wire \EXU/ALU/adder/_014_ ;
wire \EXU/ALU/adder/_015_ ;
wire \EXU/ALU/adder/_016_ ;
wire \EXU/ALU/adder/_017_ ;
wire \EXU/ALU/adder/_018_ ;
wire \EXU/ALU/adder/_019_ ;
wire \EXU/ALU/adder/_020_ ;
wire \EXU/ALU/adder/_021_ ;
wire \EXU/ALU/adder/_022_ ;
wire \EXU/ALU/adder/_023_ ;
wire \EXU/ALU/adder/_024_ ;
wire \EXU/ALU/adder/_025_ ;
wire \EXU/ALU/adder/_026_ ;
wire \EXU/ALU/adder/_027_ ;
wire \EXU/ALU/adder/_028_ ;
wire \EXU/ALU/adder/_029_ ;
wire \EXU/ALU/adder/_030_ ;
wire \EXU/ALU/adder/_031_ ;
wire \EXU/ALU/adder/_032_ ;
wire \EXU/ALU/adder/_033_ ;
wire \EXU/ALU/adder/_034_ ;
wire \EXU/ALU/adder/_035_ ;
wire \EXU/ALU/adder/_036_ ;
wire \EXU/ALU/adder/_037_ ;
wire \EXU/ALU/adder/_038_ ;
wire \EXU/ALU/adder/_039_ ;
wire \EXU/ALU/adder/_040_ ;
wire \EXU/ALU/adder/_041_ ;
wire \EXU/ALU/adder/_042_ ;
wire \EXU/ALU/adder/_043_ ;
wire \EXU/ALU/adder/_044_ ;
wire \EXU/ALU/adder/_045_ ;
wire \EXU/ALU/adder/_046_ ;
wire \EXU/ALU/adder/_047_ ;
wire \EXU/ALU/adder/_048_ ;
wire \EXU/ALU/adder/_049_ ;
wire \EXU/ALU/adder/_050_ ;
wire \EXU/ALU/adder/_051_ ;
wire \EXU/ALU/adder/_052_ ;
wire \EXU/ALU/adder/_053_ ;
wire \EXU/ALU/adder/_054_ ;
wire \EXU/ALU/adder/_055_ ;
wire \EXU/ALU/adder/_056_ ;
wire \EXU/ALU/adder/_057_ ;
wire \EXU/ALU/adder/_058_ ;
wire \EXU/ALU/adder/_059_ ;
wire \EXU/ALU/adder/_060_ ;
wire \EXU/ALU/adder/_061_ ;
wire \EXU/ALU/adder/_062_ ;
wire \EXU/ALU/adder/_063_ ;
wire \EXU/ALU/adder/_064_ ;
wire \EXU/ALU/adder/_065_ ;
wire \EXU/ALU/adder/_066_ ;
wire \EXU/ALU/adder/_067_ ;
wire \EXU/ALU/adder/_068_ ;
wire \EXU/ALU/adder/_069_ ;
wire \EXU/ALU/adder/_070_ ;
wire \EXU/ALU/adder/_071_ ;
wire \EXU/ALU/adder/_072_ ;
wire \EXU/ALU/adder/_073_ ;
wire \EXU/ALU/adder/_074_ ;
wire \EXU/ALU/adder/_075_ ;
wire \EXU/ALU/adder/_076_ ;
wire \EXU/ALU/adder/_077_ ;
wire \EXU/ALU/adder/_078_ ;
wire \EXU/ALU/adder/_079_ ;
wire \EXU/ALU/adder/_080_ ;
wire \EXU/ALU/adder/_081_ ;
wire \EXU/ALU/adder/_082_ ;
wire \EXU/ALU/adder/_083_ ;
wire \EXU/ALU/adder/_084_ ;
wire \EXU/ALU/adder/_085_ ;
wire \EXU/ALU/adder/_086_ ;
wire \EXU/ALU/adder/_087_ ;
wire \EXU/ALU/adder/_088_ ;
wire \EXU/ALU/adder/_089_ ;
wire \EXU/ALU/adder/_090_ ;
wire \EXU/ALU/adder/_091_ ;
wire \EXU/ALU/adder/_092_ ;
wire \EXU/ALU/adder/_093_ ;
wire \EXU/ALU/adder/_094_ ;
wire \EXU/ALU/adder/_095_ ;
wire \EXU/ALU/adder/_096_ ;
wire \EXU/ALU/adder/_097_ ;
wire \EXU/ALU/adder/_098_ ;
wire \EXU/ALU/adder/_099_ ;
wire \EXU/ALU/adder/_100_ ;
wire \EXU/ALU/adder/_101_ ;
wire \EXU/ALU/adder/_102_ ;
wire \EXU/ALU/adder/_103_ ;
wire \EXU/ALU/adder/_104_ ;
wire \EXU/ALU/adder/_105_ ;
wire \EXU/ALU/adder/_106_ ;
wire \EXU/ALU/adder/_107_ ;
wire \EXU/ALU/adder/_108_ ;
wire \EXU/ALU/adder/_109_ ;
wire \EXU/ALU/adder/_110_ ;
wire \EXU/ALU/adder/_111_ ;
wire \EXU/ALU/adder/_112_ ;
wire \EXU/ALU/adder/_113_ ;
wire \EXU/ALU/adder/_114_ ;
wire \EXU/ALU/adder/_115_ ;
wire \EXU/ALU/adder/_116_ ;
wire \EXU/ALU/adder/_117_ ;
wire \EXU/ALU/adder/_118_ ;
wire \EXU/ALU/adder/_119_ ;
wire \EXU/ALU/adder/_120_ ;
wire \EXU/ALU/adder/_121_ ;
wire \EXU/ALU/adder/_122_ ;
wire \EXU/ALU/adder/_123_ ;
wire \EXU/ALU/adder/_124_ ;
wire \EXU/ALU/adder/_125_ ;
wire \EXU/ALU/adder/_126_ ;
wire \EXU/ALU/adder/_127_ ;
wire \EXU/ALU/adder/_128_ ;
wire \EXU/ALU/adder/_129_ ;
wire \EXU/ALU/adder/_130_ ;
wire \EXU/ALU/adder/_131_ ;
wire \EXU/ALU/adder/_132_ ;
wire \EXU/ALU/adder/_133_ ;
wire \EXU/ALU/adder/_134_ ;
wire \EXU/ALU/adder/_135_ ;
wire \EXU/ALU/adder/_136_ ;
wire \EXU/ALU/adder/_137_ ;
wire \EXU/ALU/adder/_138_ ;
wire \EXU/ALU/adder/_139_ ;
wire \EXU/ALU/adder/_140_ ;
wire \EXU/ALU/adder/_141_ ;
wire \EXU/ALU/adder/_142_ ;
wire \EXU/ALU/adder/_143_ ;
wire \EXU/ALU/adder/_144_ ;
wire \EXU/ALU/adder/_145_ ;
wire \EXU/ALU/adder/_146_ ;
wire \EXU/ALU/adder/_147_ ;
wire \EXU/ALU/adder/_148_ ;
wire \EXU/ALU/adder/_149_ ;
wire \EXU/ALU/adder/_150_ ;
wire \EXU/ALU/adder/_151_ ;
wire \EXU/ALU/adder/_152_ ;
wire \EXU/ALU/adder/_153_ ;
wire \EXU/ALU/adder/_154_ ;
wire \EXU/ALU/adder/_155_ ;
wire \EXU/ALU/adder/_156_ ;
wire \EXU/ALU/adder/_157_ ;
wire \EXU/ALU/adder/_158_ ;
wire \EXU/ALU/adder/_159_ ;
wire \EXU/ALU/adder/_160_ ;
wire \EXU/ALU/adder/_161_ ;
wire \EXU/ALU/adder/_162_ ;
wire \EXU/ALU/adder/_163_ ;
wire \EXU/ALU/adder/_164_ ;
wire \EXU/ALU/adder/_165_ ;
wire \EXU/ALU/adder/_166_ ;
wire \EXU/ALU/adder/_167_ ;
wire \EXU/ALU/adder/_168_ ;
wire \EXU/ALU/adder/_169_ ;
wire \EXU/ALU/adder/_170_ ;
wire \EXU/ALU/adder/_171_ ;
wire \EXU/ALU/adder/_172_ ;
wire \EXU/ALU/adder/_173_ ;
wire \EXU/ALU/adder/_174_ ;
wire \EXU/ALU/adder/_175_ ;
wire \EXU/ALU/adder/_176_ ;
wire \EXU/ALU/adder/_177_ ;
wire \EXU/ALU/adder/_178_ ;
wire \EXU/ALU/adder/_179_ ;
wire \EXU/ALU/adder/_180_ ;
wire \EXU/ALU/adder/_181_ ;
wire \EXU/ALU/adder/_182_ ;
wire \EXU/ALU/adder/_183_ ;
wire \EXU/ALU/adder/_184_ ;
wire \EXU/ALU/adder/_185_ ;
wire \EXU/ALU/adder/_186_ ;
wire \EXU/ALU/adder/_187_ ;
wire \EXU/ALU/adder/_188_ ;
wire \EXU/ALU/adder/_189_ ;
wire \EXU/ALU/adder/_190_ ;
wire \EXU/ALU/adder/_191_ ;
wire \EXU/ALU/adder/_192_ ;
wire \EXU/ALU/adder/_193_ ;
wire \EXU/ALU/adder/_194_ ;
wire \EXU/ALU/adder/_195_ ;
wire \EXU/ALU/adder/_196_ ;
wire \EXU/ALU/adder/_197_ ;
wire \EXU/ALU/adder/_198_ ;
wire \EXU/ALU/adder/_199_ ;
wire \EXU/ALU/adder/_200_ ;
wire \EXU/ALU/adder/_201_ ;
wire \EXU/ALU/adder/_202_ ;
wire \EXU/ALU/adder/_203_ ;
wire \EXU/ALU/adder/_204_ ;
wire \EXU/ALU/adder/_205_ ;
wire \EXU/ALU/adder/_206_ ;
wire \EXU/ALU/adder/_207_ ;
wire \EXU/ALU/adder/_208_ ;
wire \EXU/ALU/adder/_209_ ;
wire \EXU/ALU/adder/_210_ ;
wire \EXU/ALU/adder/_211_ ;
wire \EXU/ALU/adder/_212_ ;
wire \EXU/ALU/adder/_213_ ;
wire \EXU/ALU/adder/_214_ ;
wire \EXU/ALU/adder/_215_ ;
wire \EXU/ALU/adder/_216_ ;
wire \EXU/ALU/adder/_217_ ;
wire \EXU/ALU/adder/_218_ ;
wire \EXU/ALU/adder/_219_ ;
wire \EXU/ALU/adder/_220_ ;
wire \EXU/ALU/adder/_221_ ;
wire \EXU/ALU/adder/_222_ ;
wire \EXU/ALU/adder/_223_ ;
wire \EXU/ALU/adder/_224_ ;
wire \EXU/ALU/adder/_225_ ;
wire \EXU/ALU/adder/_226_ ;
wire \EXU/ALU/adder/_227_ ;
wire \EXU/ALU/adder/_228_ ;
wire \EXU/ALU/adder/_229_ ;
wire \EXU/ALU/adder/_230_ ;
wire \EXU/ALU/adder/_231_ ;
wire \EXU/ALU/adder/_232_ ;
wire \EXU/ALU/adder/_233_ ;
wire \EXU/ALU/adder/_234_ ;
wire \EXU/ALU/adder/_235_ ;
wire \EXU/ALU/adder/_236_ ;
wire \EXU/ALU/adder/_237_ ;
wire \EXU/ALU/adder/_238_ ;
wire \EXU/ALU/adder/_239_ ;
wire \EXU/ALU/adder/_240_ ;
wire \EXU/ALU/adder/_241_ ;
wire \EXU/ALU/adder/_242_ ;
wire \EXU/ALU/adder/_243_ ;
wire \EXU/ALU/adder/_244_ ;
wire \EXU/ALU/adder/_245_ ;
wire \EXU/ALU/adder/_246_ ;
wire \EXU/ALU/adder/_247_ ;
wire \EXU/ALU/adder/_248_ ;
wire \EXU/ALU/adder/_249_ ;
wire \EXU/ALU/adder/_250_ ;
wire \EXU/ALU/adder/_251_ ;
wire \EXU/ALU/adder/_252_ ;
wire \EXU/ALU/adder/_253_ ;
wire \EXU/ALU/adder/_254_ ;
wire \EXU/ALU/adder/_255_ ;
wire \EXU/ALU/adder/_256_ ;
wire \EXU/ALU/adder/_257_ ;
wire \EXU/ALU/adder/_258_ ;
wire \EXU/ALU/adder/_259_ ;
wire \EXU/ALU/adder/_260_ ;
wire \EXU/ALU/adder/_261_ ;
wire \EXU/ALU/adder/_262_ ;
wire \EXU/ALU/adder/_263_ ;
wire \EXU/ALU/adder/_264_ ;
wire \EXU/ALU/adder/_265_ ;
wire \EXU/ALU/adder/_266_ ;
wire \EXU/ALU/adder/_267_ ;
wire \EXU/ALU/adder/_268_ ;
wire \EXU/ALU/adder/_269_ ;
wire \EXU/ALU/adder/_270_ ;
wire \EXU/ALU/adder/_271_ ;
wire \EXU/ALU/adder/_272_ ;
wire \EXU/ALU/adder/_273_ ;
wire \EXU/ALU/adder/_274_ ;
wire \EXU/ALU/adder/_275_ ;
wire \EXU/ALU/adder/_276_ ;
wire \EXU/ALU/adder/_277_ ;
wire \EXU/ALU/adder/_278_ ;
wire \EXU/ALU/adder/_279_ ;
wire \EXU/ALU/adder/_280_ ;
wire \EXU/ALU/adder/_281_ ;
wire \EXU/ALU/adder/_282_ ;
wire \EXU/ALU/adder/_283_ ;
wire \EXU/ALU/adder/_284_ ;
wire \EXU/ALU/adder/_285_ ;
wire \EXU/ALU/adder/_286_ ;
wire \EXU/ALU/adder/_287_ ;
wire \EXU/ALU/adder/_288_ ;
wire \EXU/ALU/adder/_289_ ;
wire \EXU/ALU/adder/_290_ ;
wire \EXU/ALU/adder/_291_ ;
wire \EXU/ALU/adder/_292_ ;
wire \EXU/ALU/adder/_293_ ;
wire \EXU/ALU/adder/_294_ ;
wire \EXU/ALU/adder/_295_ ;
wire \EXU/ALU/adder/_296_ ;
wire \EXU/ALU/adder/_297_ ;
wire \EXU/ALU/adder/_298_ ;
wire \EXU/ALU/adder/_299_ ;
wire \EXU/ALU/adder/_300_ ;
wire \EXU/ALU/adder/_301_ ;
wire \EXU/ALU/adder/_302_ ;
wire \EXU/ALU/adder/_303_ ;
wire \EXU/ALU/adder/_304_ ;
wire \EXU/ALU/adder/_305_ ;
wire \EXU/ALU/adder/_306_ ;
wire \EXU/ALU/adder/_307_ ;
wire \EXU/ALU/adder/_308_ ;
wire \EXU/ALU/adder/_309_ ;
wire \EXU/ALU/adder/_310_ ;
wire \EXU/ALU/adder/_311_ ;
wire \EXU/ALU/adder/_312_ ;
wire \EXU/ALU/adder/_313_ ;
wire \EXU/ALU/adder/_314_ ;
wire \EXU/ALU/adder/_315_ ;
wire \EXU/ALU/adder/_316_ ;
wire \EXU/ALU/adder/_317_ ;
wire \EXU/ALU/adder/_318_ ;
wire \EXU/ALU/adder/_319_ ;
wire \EXU/ALU/adder/_320_ ;
wire \EXU/ALU/adder/_321_ ;
wire \EXU/ALU/adder/_322_ ;
wire \EXU/ALU/adder/_323_ ;
wire \EXU/ALU/adder/_324_ ;
wire \EXU/ALU/adder/_325_ ;
wire \EXU/ALU/adder/_326_ ;
wire \EXU/ALU/adder/_327_ ;
wire \EXU/ALU/adder/_328_ ;
wire \EXU/ALU/adder/_329_ ;
wire \EXU/ALU/adder/_330_ ;
wire \EXU/ALU/adder/_331_ ;
wire \EXU/ALU/adder/_332_ ;
wire \EXU/ALU/adder/_333_ ;
wire \EXU/ALU/adder/_334_ ;
wire \EXU/ALU/adder/_335_ ;
wire \EXU/ALU/adder/_336_ ;
wire \EXU/ALU/adder/_337_ ;
wire \EXU/ALU/adder/_338_ ;
wire \EXU/ALU/adder/_339_ ;
wire \EXU/ALU/adder/_340_ ;
wire \EXU/ALU/adder/_341_ ;
wire \EXU/ALU/adder/_342_ ;
wire \EXU/ALU/adder/_343_ ;
wire \EXU/ALU/adder/_344_ ;
wire \EXU/ALU/adder/_345_ ;
wire \EXU/ALU/adder/_346_ ;
wire \EXU/ALU/adder/_347_ ;
wire \EXU/ALU/adder/_348_ ;
wire \EXU/ALU/adder/_349_ ;
wire \EXU/ALU/adder/_350_ ;
wire \EXU/ALU/adder/_351_ ;
wire \EXU/ALU/adder/_352_ ;
wire \EXU/ALU/adder/_353_ ;
wire \EXU/ALU/adder/_354_ ;
wire \EXU/ALU/adder/_355_ ;
wire \EXU/ALU/adder/_356_ ;
wire \EXU/ALU/adder/_357_ ;
wire \EXU/ALU/adder/_358_ ;
wire \EXU/ALU/adder/_359_ ;
wire \EXU/ALU/adder/_360_ ;
wire \EXU/ALU/adder/_361_ ;
wire \EXU/ALU/adder/_362_ ;
wire \EXU/ALU/adder/_363_ ;
wire \EXU/ALU/adder/_364_ ;
wire \EXU/ALU/adder/_365_ ;
wire \EXU/ALU/adder/_366_ ;
wire \EXU/ALU/adder/_367_ ;
wire \EXU/ALU/adder/_368_ ;
wire \EXU/ALU/adder/_369_ ;
wire \EXU/ALU/adder/_370_ ;
wire \EXU/ALU/aluControl/_00_ ;
wire \EXU/ALU/aluControl/_01_ ;
wire \EXU/ALU/aluControl/_02_ ;
wire \EXU/ALU/aluControl/_03_ ;
wire \EXU/ALU/aluControl/_04_ ;
wire \EXU/ALU/barrelShift/_0000_ ;
wire \EXU/ALU/barrelShift/_0001_ ;
wire \EXU/ALU/barrelShift/_0002_ ;
wire \EXU/ALU/barrelShift/_0003_ ;
wire \EXU/ALU/barrelShift/_0004_ ;
wire \EXU/ALU/barrelShift/_0005_ ;
wire \EXU/ALU/barrelShift/_0006_ ;
wire \EXU/ALU/barrelShift/_0007_ ;
wire \EXU/ALU/barrelShift/_0008_ ;
wire \EXU/ALU/barrelShift/_0009_ ;
wire \EXU/ALU/barrelShift/_0010_ ;
wire \EXU/ALU/barrelShift/_0011_ ;
wire \EXU/ALU/barrelShift/_0012_ ;
wire \EXU/ALU/barrelShift/_0013_ ;
wire \EXU/ALU/barrelShift/_0014_ ;
wire \EXU/ALU/barrelShift/_0015_ ;
wire \EXU/ALU/barrelShift/_0016_ ;
wire \EXU/ALU/barrelShift/_0017_ ;
wire \EXU/ALU/barrelShift/_0018_ ;
wire \EXU/ALU/barrelShift/_0019_ ;
wire \EXU/ALU/barrelShift/_0020_ ;
wire \EXU/ALU/barrelShift/_0021_ ;
wire \EXU/ALU/barrelShift/_0022_ ;
wire \EXU/ALU/barrelShift/_0023_ ;
wire \EXU/ALU/barrelShift/_0024_ ;
wire \EXU/ALU/barrelShift/_0025_ ;
wire \EXU/ALU/barrelShift/_0026_ ;
wire \EXU/ALU/barrelShift/_0027_ ;
wire \EXU/ALU/barrelShift/_0028_ ;
wire \EXU/ALU/barrelShift/_0029_ ;
wire \EXU/ALU/barrelShift/_0030_ ;
wire \EXU/ALU/barrelShift/_0031_ ;
wire \EXU/ALU/barrelShift/_0032_ ;
wire \EXU/ALU/barrelShift/_0033_ ;
wire \EXU/ALU/barrelShift/_0034_ ;
wire \EXU/ALU/barrelShift/_0035_ ;
wire \EXU/ALU/barrelShift/_0036_ ;
wire \EXU/ALU/barrelShift/_0037_ ;
wire \EXU/ALU/barrelShift/_0038_ ;
wire \EXU/ALU/barrelShift/_0039_ ;
wire \EXU/ALU/barrelShift/_0040_ ;
wire \EXU/ALU/barrelShift/_0041_ ;
wire \EXU/ALU/barrelShift/_0042_ ;
wire \EXU/ALU/barrelShift/_0043_ ;
wire \EXU/ALU/barrelShift/_0044_ ;
wire \EXU/ALU/barrelShift/_0045_ ;
wire \EXU/ALU/barrelShift/_0046_ ;
wire \EXU/ALU/barrelShift/_0047_ ;
wire \EXU/ALU/barrelShift/_0048_ ;
wire \EXU/ALU/barrelShift/_0049_ ;
wire \EXU/ALU/barrelShift/_0050_ ;
wire \EXU/ALU/barrelShift/_0051_ ;
wire \EXU/ALU/barrelShift/_0052_ ;
wire \EXU/ALU/barrelShift/_0053_ ;
wire \EXU/ALU/barrelShift/_0054_ ;
wire \EXU/ALU/barrelShift/_0055_ ;
wire \EXU/ALU/barrelShift/_0056_ ;
wire \EXU/ALU/barrelShift/_0057_ ;
wire \EXU/ALU/barrelShift/_0058_ ;
wire \EXU/ALU/barrelShift/_0059_ ;
wire \EXU/ALU/barrelShift/_0060_ ;
wire \EXU/ALU/barrelShift/_0061_ ;
wire \EXU/ALU/barrelShift/_0062_ ;
wire \EXU/ALU/barrelShift/_0063_ ;
wire \EXU/ALU/barrelShift/_0064_ ;
wire \EXU/ALU/barrelShift/_0065_ ;
wire \EXU/ALU/barrelShift/_0066_ ;
wire \EXU/ALU/barrelShift/_0067_ ;
wire \EXU/ALU/barrelShift/_0068_ ;
wire \EXU/ALU/barrelShift/_0069_ ;
wire \EXU/ALU/barrelShift/_0070_ ;
wire \EXU/ALU/barrelShift/_0071_ ;
wire \EXU/ALU/barrelShift/_0072_ ;
wire \EXU/ALU/barrelShift/_0073_ ;
wire \EXU/ALU/barrelShift/_0074_ ;
wire \EXU/ALU/barrelShift/_0075_ ;
wire \EXU/ALU/barrelShift/_0076_ ;
wire \EXU/ALU/barrelShift/_0077_ ;
wire \EXU/ALU/barrelShift/_0078_ ;
wire \EXU/ALU/barrelShift/_0079_ ;
wire \EXU/ALU/barrelShift/_0080_ ;
wire \EXU/ALU/barrelShift/_0081_ ;
wire \EXU/ALU/barrelShift/_0082_ ;
wire \EXU/ALU/barrelShift/_0083_ ;
wire \EXU/ALU/barrelShift/_0084_ ;
wire \EXU/ALU/barrelShift/_0085_ ;
wire \EXU/ALU/barrelShift/_0086_ ;
wire \EXU/ALU/barrelShift/_0087_ ;
wire \EXU/ALU/barrelShift/_0088_ ;
wire \EXU/ALU/barrelShift/_0089_ ;
wire \EXU/ALU/barrelShift/_0090_ ;
wire \EXU/ALU/barrelShift/_0091_ ;
wire \EXU/ALU/barrelShift/_0092_ ;
wire \EXU/ALU/barrelShift/_0093_ ;
wire \EXU/ALU/barrelShift/_0094_ ;
wire \EXU/ALU/barrelShift/_0095_ ;
wire \EXU/ALU/barrelShift/_0096_ ;
wire \EXU/ALU/barrelShift/_0097_ ;
wire \EXU/ALU/barrelShift/_0098_ ;
wire \EXU/ALU/barrelShift/_0099_ ;
wire \EXU/ALU/barrelShift/_0100_ ;
wire \EXU/ALU/barrelShift/_0101_ ;
wire \EXU/ALU/barrelShift/_0102_ ;
wire \EXU/ALU/barrelShift/_0103_ ;
wire \EXU/ALU/barrelShift/_0104_ ;
wire \EXU/ALU/barrelShift/_0105_ ;
wire \EXU/ALU/barrelShift/_0106_ ;
wire \EXU/ALU/barrelShift/_0107_ ;
wire \EXU/ALU/barrelShift/_0108_ ;
wire \EXU/ALU/barrelShift/_0109_ ;
wire \EXU/ALU/barrelShift/_0110_ ;
wire \EXU/ALU/barrelShift/_0111_ ;
wire \EXU/ALU/barrelShift/_0112_ ;
wire \EXU/ALU/barrelShift/_0113_ ;
wire \EXU/ALU/barrelShift/_0114_ ;
wire \EXU/ALU/barrelShift/_0115_ ;
wire \EXU/ALU/barrelShift/_0116_ ;
wire \EXU/ALU/barrelShift/_0117_ ;
wire \EXU/ALU/barrelShift/_0118_ ;
wire \EXU/ALU/barrelShift/_0119_ ;
wire \EXU/ALU/barrelShift/_0120_ ;
wire \EXU/ALU/barrelShift/_0121_ ;
wire \EXU/ALU/barrelShift/_0122_ ;
wire \EXU/ALU/barrelShift/_0123_ ;
wire \EXU/ALU/barrelShift/_0124_ ;
wire \EXU/ALU/barrelShift/_0125_ ;
wire \EXU/ALU/barrelShift/_0126_ ;
wire \EXU/ALU/barrelShift/_0127_ ;
wire \EXU/ALU/barrelShift/_0128_ ;
wire \EXU/ALU/barrelShift/_0129_ ;
wire \EXU/ALU/barrelShift/_0130_ ;
wire \EXU/ALU/barrelShift/_0131_ ;
wire \EXU/ALU/barrelShift/_0132_ ;
wire \EXU/ALU/barrelShift/_0133_ ;
wire \EXU/ALU/barrelShift/_0134_ ;
wire \EXU/ALU/barrelShift/_0135_ ;
wire \EXU/ALU/barrelShift/_0136_ ;
wire \EXU/ALU/barrelShift/_0137_ ;
wire \EXU/ALU/barrelShift/_0138_ ;
wire \EXU/ALU/barrelShift/_0139_ ;
wire \EXU/ALU/barrelShift/_0140_ ;
wire \EXU/ALU/barrelShift/_0141_ ;
wire \EXU/ALU/barrelShift/_0142_ ;
wire \EXU/ALU/barrelShift/_0143_ ;
wire \EXU/ALU/barrelShift/_0144_ ;
wire \EXU/ALU/barrelShift/_0145_ ;
wire \EXU/ALU/barrelShift/_0146_ ;
wire \EXU/ALU/barrelShift/_0147_ ;
wire \EXU/ALU/barrelShift/_0148_ ;
wire \EXU/ALU/barrelShift/_0149_ ;
wire \EXU/ALU/barrelShift/_0150_ ;
wire \EXU/ALU/barrelShift/_0151_ ;
wire \EXU/ALU/barrelShift/_0152_ ;
wire \EXU/ALU/barrelShift/_0153_ ;
wire \EXU/ALU/barrelShift/_0154_ ;
wire \EXU/ALU/barrelShift/_0155_ ;
wire \EXU/ALU/barrelShift/_0156_ ;
wire \EXU/ALU/barrelShift/_0157_ ;
wire \EXU/ALU/barrelShift/_0158_ ;
wire \EXU/ALU/barrelShift/_0159_ ;
wire \EXU/ALU/barrelShift/_0160_ ;
wire \EXU/ALU/barrelShift/_0161_ ;
wire \EXU/ALU/barrelShift/_0162_ ;
wire \EXU/ALU/barrelShift/_0163_ ;
wire \EXU/ALU/barrelShift/_0164_ ;
wire \EXU/ALU/barrelShift/_0165_ ;
wire \EXU/ALU/barrelShift/_0166_ ;
wire \EXU/ALU/barrelShift/_0167_ ;
wire \EXU/ALU/barrelShift/_0168_ ;
wire \EXU/ALU/barrelShift/_0169_ ;
wire \EXU/ALU/barrelShift/_0170_ ;
wire \EXU/ALU/barrelShift/_0171_ ;
wire \EXU/ALU/barrelShift/_0172_ ;
wire \EXU/ALU/barrelShift/_0173_ ;
wire \EXU/ALU/barrelShift/_0174_ ;
wire \EXU/ALU/barrelShift/_0175_ ;
wire \EXU/ALU/barrelShift/_0176_ ;
wire \EXU/ALU/barrelShift/_0177_ ;
wire \EXU/ALU/barrelShift/_0178_ ;
wire \EXU/ALU/barrelShift/_0179_ ;
wire \EXU/ALU/barrelShift/_0180_ ;
wire \EXU/ALU/barrelShift/_0181_ ;
wire \EXU/ALU/barrelShift/_0182_ ;
wire \EXU/ALU/barrelShift/_0183_ ;
wire \EXU/ALU/barrelShift/_0184_ ;
wire \EXU/ALU/barrelShift/_0185_ ;
wire \EXU/ALU/barrelShift/_0186_ ;
wire \EXU/ALU/barrelShift/_0187_ ;
wire \EXU/ALU/barrelShift/_0188_ ;
wire \EXU/ALU/barrelShift/_0189_ ;
wire \EXU/ALU/barrelShift/_0190_ ;
wire \EXU/ALU/barrelShift/_0191_ ;
wire \EXU/ALU/barrelShift/_0192_ ;
wire \EXU/ALU/barrelShift/_0193_ ;
wire \EXU/ALU/barrelShift/_0194_ ;
wire \EXU/ALU/barrelShift/_0195_ ;
wire \EXU/ALU/barrelShift/_0196_ ;
wire \EXU/ALU/barrelShift/_0197_ ;
wire \EXU/ALU/barrelShift/_0198_ ;
wire \EXU/ALU/barrelShift/_0199_ ;
wire \EXU/ALU/barrelShift/_0200_ ;
wire \EXU/ALU/barrelShift/_0201_ ;
wire \EXU/ALU/barrelShift/_0202_ ;
wire \EXU/ALU/barrelShift/_0203_ ;
wire \EXU/ALU/barrelShift/_0204_ ;
wire \EXU/ALU/barrelShift/_0205_ ;
wire \EXU/ALU/barrelShift/_0206_ ;
wire \EXU/ALU/barrelShift/_0207_ ;
wire \EXU/ALU/barrelShift/_0208_ ;
wire \EXU/ALU/barrelShift/_0209_ ;
wire \EXU/ALU/barrelShift/_0210_ ;
wire \EXU/ALU/barrelShift/_0211_ ;
wire \EXU/ALU/barrelShift/_0212_ ;
wire \EXU/ALU/barrelShift/_0213_ ;
wire \EXU/ALU/barrelShift/_0214_ ;
wire \EXU/ALU/barrelShift/_0215_ ;
wire \EXU/ALU/barrelShift/_0216_ ;
wire \EXU/ALU/barrelShift/_0217_ ;
wire \EXU/ALU/barrelShift/_0218_ ;
wire \EXU/ALU/barrelShift/_0219_ ;
wire \EXU/ALU/barrelShift/_0220_ ;
wire \EXU/ALU/barrelShift/_0221_ ;
wire \EXU/ALU/barrelShift/_0222_ ;
wire \EXU/ALU/barrelShift/_0223_ ;
wire \EXU/ALU/barrelShift/_0224_ ;
wire \EXU/ALU/barrelShift/_0225_ ;
wire \EXU/ALU/barrelShift/_0226_ ;
wire \EXU/ALU/barrelShift/_0227_ ;
wire \EXU/ALU/barrelShift/_0228_ ;
wire \EXU/ALU/barrelShift/_0229_ ;
wire \EXU/ALU/barrelShift/_0230_ ;
wire \EXU/ALU/barrelShift/_0231_ ;
wire \EXU/ALU/barrelShift/_0232_ ;
wire \EXU/ALU/barrelShift/_0233_ ;
wire \EXU/ALU/barrelShift/_0234_ ;
wire \EXU/ALU/barrelShift/_0235_ ;
wire \EXU/ALU/barrelShift/_0236_ ;
wire \EXU/ALU/barrelShift/_0237_ ;
wire \EXU/ALU/barrelShift/_0238_ ;
wire \EXU/ALU/barrelShift/_0239_ ;
wire \EXU/ALU/barrelShift/_0240_ ;
wire \EXU/ALU/barrelShift/_0241_ ;
wire \EXU/ALU/barrelShift/_0242_ ;
wire \EXU/ALU/barrelShift/_0243_ ;
wire \EXU/ALU/barrelShift/_0244_ ;
wire \EXU/ALU/barrelShift/_0245_ ;
wire \EXU/ALU/barrelShift/_0246_ ;
wire \EXU/ALU/barrelShift/_0247_ ;
wire \EXU/ALU/barrelShift/_0248_ ;
wire \EXU/ALU/barrelShift/_0249_ ;
wire \EXU/ALU/barrelShift/_0250_ ;
wire \EXU/ALU/barrelShift/_0251_ ;
wire \EXU/ALU/barrelShift/_0252_ ;
wire \EXU/ALU/barrelShift/_0253_ ;
wire \EXU/ALU/barrelShift/_0254_ ;
wire \EXU/ALU/barrelShift/_0255_ ;
wire \EXU/ALU/barrelShift/_0256_ ;
wire \EXU/ALU/barrelShift/_0257_ ;
wire \EXU/ALU/barrelShift/_0258_ ;
wire \EXU/ALU/barrelShift/_0259_ ;
wire \EXU/ALU/barrelShift/_0260_ ;
wire \EXU/ALU/barrelShift/_0261_ ;
wire \EXU/ALU/barrelShift/_0262_ ;
wire \EXU/ALU/barrelShift/_0263_ ;
wire \EXU/ALU/barrelShift/_0264_ ;
wire \EXU/ALU/barrelShift/_0265_ ;
wire \EXU/ALU/barrelShift/_0266_ ;
wire \EXU/ALU/barrelShift/_0267_ ;
wire \EXU/ALU/barrelShift/_0268_ ;
wire \EXU/ALU/barrelShift/_0269_ ;
wire \EXU/ALU/barrelShift/_0270_ ;
wire \EXU/ALU/barrelShift/_0271_ ;
wire \EXU/ALU/barrelShift/_0272_ ;
wire \EXU/ALU/barrelShift/_0273_ ;
wire \EXU/ALU/barrelShift/_0274_ ;
wire \EXU/ALU/barrelShift/_0275_ ;
wire \EXU/ALU/barrelShift/_0276_ ;
wire \EXU/ALU/barrelShift/_0277_ ;
wire \EXU/ALU/barrelShift/_0278_ ;
wire \EXU/ALU/barrelShift/_0279_ ;
wire \EXU/ALU/barrelShift/_0280_ ;
wire \EXU/ALU/barrelShift/_0281_ ;
wire \EXU/ALU/barrelShift/_0282_ ;
wire \EXU/ALU/barrelShift/_0283_ ;
wire \EXU/ALU/barrelShift/_0284_ ;
wire \EXU/ALU/barrelShift/_0285_ ;
wire \EXU/ALU/barrelShift/_0286_ ;
wire \EXU/ALU/barrelShift/_0287_ ;
wire \EXU/ALU/barrelShift/_0288_ ;
wire \EXU/ALU/barrelShift/_0289_ ;
wire \EXU/ALU/barrelShift/_0290_ ;
wire \EXU/ALU/barrelShift/_0291_ ;
wire \EXU/ALU/barrelShift/_0292_ ;
wire \EXU/ALU/barrelShift/_0293_ ;
wire \EXU/ALU/barrelShift/_0294_ ;
wire \EXU/ALU/barrelShift/_0295_ ;
wire \EXU/ALU/barrelShift/_0296_ ;
wire \EXU/ALU/barrelShift/_0297_ ;
wire \EXU/ALU/barrelShift/_0298_ ;
wire \EXU/ALU/barrelShift/_0299_ ;
wire \EXU/ALU/barrelShift/_0300_ ;
wire \EXU/ALU/barrelShift/_0301_ ;
wire \EXU/ALU/barrelShift/_0302_ ;
wire \EXU/ALU/barrelShift/_0303_ ;
wire \EXU/ALU/barrelShift/_0304_ ;
wire \EXU/ALU/barrelShift/_0305_ ;
wire \EXU/ALU/barrelShift/_0306_ ;
wire \EXU/ALU/barrelShift/_0307_ ;
wire \EXU/ALU/barrelShift/_0308_ ;
wire \EXU/ALU/barrelShift/_0309_ ;
wire \EXU/ALU/barrelShift/_0310_ ;
wire \EXU/ALU/barrelShift/_0311_ ;
wire \EXU/ALU/barrelShift/_0312_ ;
wire \EXU/ALU/barrelShift/_0313_ ;
wire \EXU/ALU/barrelShift/_0314_ ;
wire \EXU/ALU/barrelShift/_0315_ ;
wire \EXU/ALU/barrelShift/_0316_ ;
wire \EXU/ALU/barrelShift/_0317_ ;
wire \EXU/ALU/barrelShift/_0318_ ;
wire \EXU/ALU/barrelShift/_0319_ ;
wire \EXU/ALU/barrelShift/_0320_ ;
wire \EXU/ALU/barrelShift/_0321_ ;
wire \EXU/ALU/barrelShift/_0322_ ;
wire \EXU/ALU/barrelShift/_0323_ ;
wire \EXU/ALU/barrelShift/_0324_ ;
wire \EXU/ALU/barrelShift/_0325_ ;
wire \EXU/ALU/barrelShift/_0326_ ;
wire \EXU/ALU/barrelShift/_0327_ ;
wire \EXU/ALU/barrelShift/_0328_ ;
wire \EXU/ALU/barrelShift/_0329_ ;
wire \EXU/ALU/barrelShift/_0330_ ;
wire \EXU/ALU/barrelShift/_0331_ ;
wire \EXU/ALU/barrelShift/_0332_ ;
wire \EXU/ALU/barrelShift/_0333_ ;
wire \EXU/ALU/barrelShift/_0334_ ;
wire \EXU/ALU/barrelShift/_0335_ ;
wire \EXU/ALU/barrelShift/_0336_ ;
wire \EXU/ALU/barrelShift/_0337_ ;
wire \EXU/ALU/barrelShift/_0338_ ;
wire \EXU/ALU/barrelShift/_0339_ ;
wire \EXU/ALU/barrelShift/_0340_ ;
wire \EXU/ALU/barrelShift/_0341_ ;
wire \EXU/ALU/barrelShift/_0342_ ;
wire \EXU/ALU/barrelShift/_0343_ ;
wire \EXU/ALU/barrelShift/_0344_ ;
wire \EXU/ALU/barrelShift/_0345_ ;
wire \EXU/ALU/barrelShift/_0346_ ;
wire \EXU/ALU/barrelShift/_0347_ ;
wire \EXU/ALU/barrelShift/_0348_ ;
wire \EXU/ALU/barrelShift/_0349_ ;
wire \EXU/ALU/barrelShift/_0350_ ;
wire \EXU/ALU/barrelShift/_0351_ ;
wire \EXU/ALU/barrelShift/_0352_ ;
wire \EXU/ALU/barrelShift/_0353_ ;
wire \EXU/ALU/barrelShift/_0354_ ;
wire \EXU/ALU/barrelShift/_0355_ ;
wire \EXU/ALU/barrelShift/_0356_ ;
wire \EXU/ALU/barrelShift/_0357_ ;
wire \EXU/ALU/barrelShift/_0358_ ;
wire \EXU/ALU/barrelShift/_0359_ ;
wire \EXU/ALU/barrelShift/_0360_ ;
wire \EXU/ALU/barrelShift/_0361_ ;
wire \EXU/ALU/barrelShift/_0362_ ;
wire \EXU/ALU/barrelShift/_0363_ ;
wire \EXU/ALU/barrelShift/_0364_ ;
wire \EXU/ALU/barrelShift/_0365_ ;
wire \EXU/ALU/barrelShift/_0366_ ;
wire \EXU/ALU/barrelShift/_0367_ ;
wire \EXU/ALU/barrelShift/_0368_ ;
wire \EXU/ALU/barrelShift/_0369_ ;
wire \EXU/ALU/barrelShift/_0370_ ;
wire \EXU/ALU/barrelShift/_0371_ ;
wire \EXU/ALU/barrelShift/_0372_ ;
wire \EXU/ALU/barrelShift/_0373_ ;
wire \EXU/ALU/barrelShift/_0374_ ;
wire \EXU/ALU/barrelShift/_0375_ ;
wire \EXU/ALU/barrelShift/_0376_ ;
wire \EXU/ALU/barrelShift/_0377_ ;
wire \EXU/ALU/barrelShift/_0378_ ;
wire \EXU/ALU/barrelShift/_0379_ ;
wire \EXU/ALU/barrelShift/_0380_ ;
wire \EXU/ALU/barrelShift/_0381_ ;
wire \EXU/ALU/barrelShift/_0382_ ;
wire \EXU/ALU/barrelShift/_0383_ ;
wire \EXU/ALU/barrelShift/_0384_ ;
wire \EXU/ALU/barrelShift/_0385_ ;
wire \EXU/ALU/barrelShift/_0386_ ;
wire \EXU/ALU/barrelShift/_0387_ ;
wire \EXU/ALU/barrelShift/_0388_ ;
wire \EXU/ALU/barrelShift/_0389_ ;
wire \EXU/ALU/barrelShift/_0390_ ;
wire \EXU/ALU/barrelShift/_0391_ ;
wire \EXU/ALU/barrelShift/_0392_ ;
wire \EXU/ALU/barrelShift/_0393_ ;
wire \EXU/ALU/barrelShift/_0394_ ;
wire \EXU/ALU/barrelShift/_0395_ ;
wire \EXU/ALU/barrelShift/_0396_ ;
wire \EXU/ALU/barrelShift/_0397_ ;
wire \EXU/ALU/barrelShift/_0398_ ;
wire \EXU/ALU/barrelShift/_0399_ ;
wire \EXU/ALU/barrelShift/_0400_ ;
wire \EXU/ALU/barrelShift/_0401_ ;
wire \EXU/ALU/barrelShift/_0402_ ;
wire \EXU/ALU/barrelShift/_0403_ ;
wire \EXU/ALU/barrelShift/_0404_ ;
wire \EXU/ALU/barrelShift/_0405_ ;
wire \EXU/ALU/barrelShift/_0406_ ;
wire \EXU/ALU/barrelShift/_0407_ ;
wire \EXU/ALU/barrelShift/_0408_ ;
wire \EXU/ALU/barrelShift/_0409_ ;
wire \EXU/ALU/barrelShift/_0410_ ;
wire \EXU/ALU/barrelShift/_0411_ ;
wire \EXU/ALU/barrelShift/_0412_ ;
wire \EXU/ALU/barrelShift/_0413_ ;
wire \EXU/ALU/barrelShift/_0414_ ;
wire \EXU/ALU/barrelShift/_0415_ ;
wire \EXU/ALU/barrelShift/_0416_ ;
wire \EXU/ALU/barrelShift/_0417_ ;
wire \EXU/ALU/barrelShift/_0418_ ;
wire \EXU/ALU/barrelShift/_0419_ ;
wire \EXU/ALU/barrelShift/_0420_ ;
wire \EXU/ALU/barrelShift/_0421_ ;
wire \EXU/ALU/barrelShift/_0422_ ;
wire \EXU/ALU/barrelShift/_0423_ ;
wire \EXU/ALU/barrelShift/_0424_ ;
wire \EXU/ALU/barrelShift/_0425_ ;
wire \EXU/ALU/barrelShift/_0426_ ;
wire \EXU/ALU/barrelShift/_0427_ ;
wire \EXU/ALU/barrelShift/_0428_ ;
wire \EXU/ALU/barrelShift/_0429_ ;
wire \EXU/ALU/barrelShift/_0430_ ;
wire \EXU/ALU/barrelShift/_0431_ ;
wire \EXU/ALU/barrelShift/_0432_ ;
wire \EXU/ALU/barrelShift/_0433_ ;
wire \EXU/ALU/barrelShift/_0434_ ;
wire \EXU/ALU/barrelShift/_0435_ ;
wire \EXU/ALU/barrelShift/_0436_ ;
wire \EXU/ALU/barrelShift/_0437_ ;
wire \EXU/ALU/barrelShift/_0438_ ;
wire \EXU/ALU/barrelShift/_0439_ ;
wire \EXU/ALU/barrelShift/_0440_ ;
wire \EXU/ALU/barrelShift/_0441_ ;
wire \EXU/ALU/barrelShift/_0442_ ;
wire \EXU/ALU/barrelShift/_0443_ ;
wire \EXU/ALU/barrelShift/_0444_ ;
wire \EXU/ALU/barrelShift/_0445_ ;
wire \EXU/ALU/barrelShift/_0446_ ;
wire \EXU/ALU/barrelShift/_0447_ ;
wire \EXU/ALU/barrelShift/_0448_ ;
wire \EXU/ALU/barrelShift/_0449_ ;
wire \EXU/ALU/barrelShift/_0450_ ;
wire \EXU/ALU/barrelShift/_0451_ ;
wire \EXU/ALU/barrelShift/_0452_ ;
wire \EXU/ALU/barrelShift/_0453_ ;
wire \EXU/ALU/barrelShift/_0454_ ;
wire \EXU/ALU/barrelShift/_0455_ ;
wire \EXU/ALU/barrelShift/_0456_ ;
wire \EXU/ALU/barrelShift/_0457_ ;
wire \EXU/ALU/barrelShift/_0458_ ;
wire \EXU/ALU/barrelShift/_0459_ ;
wire \EXU/ALU/barrelShift/_0460_ ;
wire \EXU/ALU/barrelShift/_0461_ ;
wire \EXU/ALU/barrelShift/_0462_ ;
wire \EXU/ALU/barrelShift/_0463_ ;
wire \EXU/ALU/barrelShift/_0464_ ;
wire \EXU/ALU/barrelShift/_0465_ ;
wire \EXU/ALU/barrelShift/_0466_ ;
wire \EXU/ALU/barrelShift/_0467_ ;
wire \EXU/ALU/barrelShift/_0468_ ;
wire \EXU/ALU/barrelShift/_0469_ ;
wire \EXU/ALU/barrelShift/_0470_ ;
wire \EXU/ALU/barrelShift/_0471_ ;
wire \EXU/ALU/barrelShift/_0472_ ;
wire \EXU/ALU/barrelShift/_0473_ ;
wire \EXU/ALU/barrelShift/_0474_ ;
wire \EXU/ALU/barrelShift/_0475_ ;
wire \EXU/ALU/barrelShift/_0476_ ;
wire \EXU/ALU/barrelShift/_0477_ ;
wire \EXU/ALU/barrelShift/_0478_ ;
wire \EXU/ALU/barrelShift/_0479_ ;
wire \EXU/ALU/barrelShift/_0480_ ;
wire \EXU/ALU/barrelShift/_0481_ ;
wire \EXU/ALU/barrelShift/_0482_ ;
wire \EXU/ALU/barrelShift/_0483_ ;
wire \EXU/ALU/barrelShift/_0484_ ;
wire \EXU/ALU/barrelShift/_0485_ ;
wire \EXU/ALU/barrelShift/_0486_ ;
wire \EXU/ALU/barrelShift/_0487_ ;
wire \EXU/ALU/barrelShift/_0488_ ;
wire \EXU/ALU/barrelShift/_0489_ ;
wire \EXU/ALU/barrelShift/_0490_ ;
wire \EXU/ALU/barrelShift/_0491_ ;
wire \EXU/ALU/barrelShift/_0492_ ;
wire \EXU/ALU/barrelShift/_0493_ ;
wire \EXU/ALU/barrelShift/_0494_ ;
wire \EXU/ALU/barrelShift/_0495_ ;
wire \EXU/ALU/barrelShift/_0496_ ;
wire \EXU/ALU/barrelShift/_0497_ ;
wire \EXU/ALU/barrelShift/_0498_ ;
wire \EXU/ALU/barrelShift/_0499_ ;
wire \EXU/ALU/barrelShift/_0500_ ;
wire \EXU/ALU/barrelShift/_0501_ ;
wire \EXU/ALU/barrelShift/_0502_ ;
wire \EXU/ALU/barrelShift/_0503_ ;
wire \EXU/ALU/barrelShift/_0504_ ;
wire \EXU/ALU/barrelShift/_0505_ ;
wire \EXU/ALU/barrelShift/_0506_ ;
wire \EXU/ALU/barrelShift/_0507_ ;
wire \EXU/ALU/barrelShift/_0508_ ;
wire \EXU/ALU/barrelShift/_0509_ ;
wire \EXU/ALU/barrelShift/_0510_ ;
wire \EXU/ALU/barrelShift/_0511_ ;
wire \EXU/ALU/barrelShift/_0512_ ;
wire \EXU/ALU/barrelShift/_0513_ ;
wire \EXU/ALU/barrelShift/_0514_ ;
wire \EXU/ALU/barrelShift/_0515_ ;
wire \EXU/ALU/barrelShift/_0516_ ;
wire \EXU/ALU/barrelShift/_0517_ ;
wire \EXU/ALU/barrelShift/_0518_ ;
wire \EXU/ALU/barrelShift/_0519_ ;
wire \EXU/ALU/barrelShift/_0520_ ;
wire \EXU/ALU/barrelShift/_0521_ ;
wire \EXU/ALU/barrelShift/_0522_ ;
wire \EXU/ALU/barrelShift/_0523_ ;
wire \EXU/ALU/barrelShift/_0524_ ;
wire \EXU/ALU/barrelShift/_0525_ ;
wire \EXU/ALU/barrelShift/_0526_ ;
wire \EXU/ALU/barrelShift/_0527_ ;
wire \EXU/ALU/barrelShift/_0528_ ;
wire \EXU/ALU/barrelShift/_0529_ ;
wire \EXU/ALU/barrelShift/_0530_ ;
wire \EXU/ALU/barrelShift/_0531_ ;
wire \EXU/ALU/barrelShift/_0532_ ;
wire \EXU/ALU/barrelShift/_0533_ ;
wire \EXU/ALU/barrelShift/_0534_ ;
wire \EXU/ALU/barrelShift/_0535_ ;
wire \EXU/ALU/barrelShift/_0536_ ;
wire \EXU/ALU/barrelShift/_0537_ ;
wire \EXU/ALU/barrelShift/_0538_ ;
wire \EXU/ALU/barrelShift/_0539_ ;
wire \EXU/ALU/barrelShift/_0540_ ;
wire \EXU/ALU/barrelShift/_0541_ ;
wire \EXU/ALU/barrelShift/_0542_ ;
wire \EXU/ALU/barrelShift/_0543_ ;
wire \EXU/ALU/barrelShift/_0544_ ;
wire \EXU/ALU/barrelShift/_0545_ ;
wire \EXU/ALU/barrelShift/_0546_ ;
wire \EXU/ALU/barrelShift/_0547_ ;
wire \EXU/ALU/barrelShift/_0548_ ;
wire \EXU/ALU/barrelShift/_0549_ ;
wire \EXU/ALU/barrelShift/_0550_ ;
wire \EXU/ALU/barrelShift/_0551_ ;
wire \EXU/ALU/barrelShift/_0552_ ;
wire \EXU/ALU/barrelShift/_0553_ ;
wire \EXU/ALU/barrelShift/_0554_ ;
wire \EXU/ALU/barrelShift/_0555_ ;
wire \EXU/ALU/barrelShift/_0556_ ;
wire \EXU/ALU/barrelShift/_0557_ ;
wire \EXU/ALU/barrelShift/_0558_ ;
wire \EXU/ALU/barrelShift/_0559_ ;
wire \EXU/ALU/barrelShift/_0560_ ;
wire \EXU/ALU/barrelShift/_0561_ ;
wire \EXU/ALU/barrelShift/_0562_ ;
wire \EXU/ALU/barrelShift/_0563_ ;
wire \EXU/ALU/barrelShift/casez_tmp_127 ;
wire \EXU/ALU/barrelShift/casez_tmp_128 ;
wire \EXU/ALU/barrelShift/casez_tmp_129 ;
wire \EXU/ALU/barrelShift/casez_tmp_130 ;
wire \EXU/ALU/barrelShift/casez_tmp_131 ;
wire \EXU/ALU/barrelShift/casez_tmp_132 ;
wire \EXU/ALU/barrelShift/casez_tmp_133 ;
wire \EXU/ALU/barrelShift/casez_tmp_134 ;
wire \EXU/ALU/barrelShift/casez_tmp_135 ;
wire \EXU/ALU/barrelShift/casez_tmp_136 ;
wire \EXU/ALU/barrelShift/casez_tmp_137 ;
wire \EXU/ALU/barrelShift/casez_tmp_138 ;
wire \EXU/ALU/barrelShift/casez_tmp_139 ;
wire \EXU/ALU/barrelShift/casez_tmp_140 ;
wire \EXU/ALU/barrelShift/casez_tmp_141 ;
wire \EXU/ALU/barrelShift/casez_tmp_142 ;
wire \EXU/ALU/barrelShift/casez_tmp_143 ;
wire \EXU/ALU/barrelShift/casez_tmp_144 ;
wire \EXU/ALU/barrelShift/casez_tmp_145 ;
wire \EXU/ALU/barrelShift/casez_tmp_146 ;
wire \EXU/ALU/barrelShift/casez_tmp_147 ;
wire \EXU/ALU/barrelShift/casez_tmp_148 ;
wire \EXU/ALU/barrelShift/casez_tmp_149 ;
wire \EXU/ALU/barrelShift/casez_tmp_150 ;
wire \EXU/ALU/barrelShift/casez_tmp_151 ;
wire \EXU/ALU/barrelShift/casez_tmp_152 ;
wire \EXU/ALU/barrelShift/casez_tmp_153 ;
wire \EXU/ALU/barrelShift/casez_tmp_154 ;
wire \EXU/ALU/barrelShift/casez_tmp_155 ;
wire \EXU/ALU/barrelShift/casez_tmp_156 ;
wire \EXU/ALU/barrelShift/casez_tmp_157 ;
wire \EXU/ALU/barrelShift/casez_tmp_158 ;
wire \EXU/BrCond/_00_ ;
wire \EXU/BrCond/_01_ ;
wire \EXU/BrCond/_02_ ;
wire \EXU/BrCond/_03_ ;
wire \EXU/BrCond/_04_ ;
wire \EXU/BrCond/_05_ ;
wire \EXU/BrCond/_06_ ;
wire \EXU/BrCond/_07_ ;
wire \EXU/BrCond/_08_ ;
wire \EXU/BrCond/_09_ ;
wire \EXU/BrCond/_10_ ;
wire \EXU/BrCond/_11_ ;
wire \EXU/BrCond/_12_ ;
wire \EXU/BrCond/_13_ ;
wire \EXU/BrCond/_14_ ;
wire \EXU/BrCond/_15_ ;
wire \EXU/BrCond/_16_ ;
wire \EXU/CSRControl/_0000_ ;
wire \EXU/CSRControl/_0001_ ;
wire \EXU/CSRControl/_0002_ ;
wire \EXU/CSRControl/_0003_ ;
wire \EXU/CSRControl/_0004_ ;
wire \EXU/CSRControl/_0005_ ;
wire \EXU/CSRControl/_0006_ ;
wire \EXU/CSRControl/_0007_ ;
wire \EXU/CSRControl/_0008_ ;
wire \EXU/CSRControl/_0009_ ;
wire \EXU/CSRControl/_0010_ ;
wire \EXU/CSRControl/_0011_ ;
wire \EXU/CSRControl/_0012_ ;
wire \EXU/CSRControl/_0013_ ;
wire \EXU/CSRControl/_0014_ ;
wire \EXU/CSRControl/_0015_ ;
wire \EXU/CSRControl/_0016_ ;
wire \EXU/CSRControl/_0017_ ;
wire \EXU/CSRControl/_0018_ ;
wire \EXU/CSRControl/_0019_ ;
wire \EXU/CSRControl/_0020_ ;
wire \EXU/CSRControl/_0021_ ;
wire \EXU/CSRControl/_0022_ ;
wire \EXU/CSRControl/_0023_ ;
wire \EXU/CSRControl/_0024_ ;
wire \EXU/CSRControl/_0025_ ;
wire \EXU/CSRControl/_0026_ ;
wire \EXU/CSRControl/_0027_ ;
wire \EXU/CSRControl/_0028_ ;
wire \EXU/CSRControl/_0029_ ;
wire \EXU/CSRControl/_0030_ ;
wire \EXU/CSRControl/_0031_ ;
wire \EXU/CSRControl/_0032_ ;
wire \EXU/CSRControl/_0033_ ;
wire \EXU/CSRControl/_0034_ ;
wire \EXU/CSRControl/_0035_ ;
wire \EXU/CSRControl/_0036_ ;
wire \EXU/CSRControl/_0037_ ;
wire \EXU/CSRControl/_0038_ ;
wire \EXU/CSRControl/_0039_ ;
wire \EXU/CSRControl/_0040_ ;
wire \EXU/CSRControl/_0041_ ;
wire \EXU/CSRControl/_0042_ ;
wire \EXU/CSRControl/_0043_ ;
wire \EXU/CSRControl/_0044_ ;
wire \EXU/CSRControl/_0045_ ;
wire \EXU/CSRControl/_0046_ ;
wire \EXU/CSRControl/_0047_ ;
wire \EXU/CSRControl/_0048_ ;
wire \EXU/CSRControl/_0049_ ;
wire \EXU/CSRControl/_0050_ ;
wire \EXU/CSRControl/_0051_ ;
wire \EXU/CSRControl/_0052_ ;
wire \EXU/CSRControl/_0053_ ;
wire \EXU/CSRControl/_0054_ ;
wire \EXU/CSRControl/_0055_ ;
wire \EXU/CSRControl/_0056_ ;
wire \EXU/CSRControl/_0057_ ;
wire \EXU/CSRControl/_0058_ ;
wire \EXU/CSRControl/_0059_ ;
wire \EXU/CSRControl/_0060_ ;
wire \EXU/CSRControl/_0061_ ;
wire \EXU/CSRControl/_0062_ ;
wire \EXU/CSRControl/_0063_ ;
wire \EXU/CSRControl/_0064_ ;
wire \EXU/CSRControl/_0065_ ;
wire \EXU/CSRControl/_0066_ ;
wire \EXU/CSRControl/_0067_ ;
wire \EXU/CSRControl/_0068_ ;
wire \EXU/CSRControl/_0069_ ;
wire \EXU/CSRControl/_0070_ ;
wire \EXU/CSRControl/_0071_ ;
wire \EXU/CSRControl/_0072_ ;
wire \EXU/CSRControl/_0073_ ;
wire \EXU/CSRControl/_0074_ ;
wire \EXU/CSRControl/_0075_ ;
wire \EXU/CSRControl/_0076_ ;
wire \EXU/CSRControl/_0077_ ;
wire \EXU/CSRControl/_0078_ ;
wire \EXU/CSRControl/_0079_ ;
wire \EXU/CSRControl/_0080_ ;
wire \EXU/CSRControl/_0081_ ;
wire \EXU/CSRControl/_0082_ ;
wire \EXU/CSRControl/_0083_ ;
wire \EXU/CSRControl/_0084_ ;
wire \EXU/CSRControl/_0085_ ;
wire \EXU/CSRControl/_0086_ ;
wire \EXU/CSRControl/_0087_ ;
wire \EXU/CSRControl/_0088_ ;
wire \EXU/CSRControl/_0089_ ;
wire \EXU/CSRControl/_0090_ ;
wire \EXU/CSRControl/_0091_ ;
wire \EXU/CSRControl/_0092_ ;
wire \EXU/CSRControl/_0093_ ;
wire \EXU/CSRControl/_0094_ ;
wire \EXU/CSRControl/_0095_ ;
wire \EXU/CSRControl/_0096_ ;
wire \EXU/CSRControl/_0097_ ;
wire \EXU/CSRControl/_0098_ ;
wire \EXU/CSRControl/_0099_ ;
wire \EXU/CSRControl/_0100_ ;
wire \EXU/CSRControl/_0101_ ;
wire \EXU/CSRControl/_0102_ ;
wire \EXU/CSRControl/_0103_ ;
wire \EXU/CSRControl/_0104_ ;
wire \EXU/CSRControl/_0105_ ;
wire \EXU/CSRControl/_0106_ ;
wire \EXU/CSRControl/_0107_ ;
wire \EXU/CSRControl/_0108_ ;
wire \EXU/CSRControl/_0109_ ;
wire \EXU/CSRControl/_0110_ ;
wire \EXU/CSRControl/_0111_ ;
wire \EXU/CSRControl/_0112_ ;
wire \EXU/CSRControl/_0113_ ;
wire \EXU/CSRControl/_0114_ ;
wire \EXU/CSRControl/_0115_ ;
wire \EXU/CSRControl/_0116_ ;
wire \EXU/CSRControl/_0117_ ;
wire \EXU/CSRControl/_0118_ ;
wire \EXU/CSRControl/_0119_ ;
wire \EXU/CSRControl/_0120_ ;
wire \EXU/CSRControl/_0121_ ;
wire \EXU/CSRControl/_0122_ ;
wire \EXU/CSRControl/_0123_ ;
wire \EXU/CSRControl/_0124_ ;
wire \EXU/CSRControl/_0125_ ;
wire \EXU/CSRControl/_0126_ ;
wire \EXU/CSRControl/_0127_ ;
wire \EXU/CSRControl/_0128_ ;
wire \EXU/CSRControl/_0129_ ;
wire \EXU/CSRControl/_0130_ ;
wire \EXU/CSRControl/_0131_ ;
wire \EXU/CSRControl/_0132_ ;
wire \EXU/CSRControl/_0133_ ;
wire \EXU/CSRControl/_0134_ ;
wire \EXU/CSRControl/_0135_ ;
wire \EXU/CSRControl/_0136_ ;
wire \EXU/CSRControl/_0137_ ;
wire \EXU/CSRControl/_0138_ ;
wire \EXU/CSRControl/_0139_ ;
wire \EXU/CSRControl/_0140_ ;
wire \EXU/CSRControl/_0141_ ;
wire \EXU/CSRControl/_0142_ ;
wire \EXU/CSRControl/_0143_ ;
wire \EXU/CSRControl/_0144_ ;
wire \EXU/CSRControl/_0145_ ;
wire \EXU/CSRControl/_0146_ ;
wire \EXU/CSRControl/_0147_ ;
wire \EXU/CSRControl/_0148_ ;
wire \EXU/CSRControl/_0149_ ;
wire \EXU/CSRControl/_0150_ ;
wire \EXU/CSRControl/_0151_ ;
wire \EXU/CSRControl/_0152_ ;
wire \EXU/CSRControl/_0153_ ;
wire \EXU/CSRControl/_0154_ ;
wire \EXU/CSRControl/_0155_ ;
wire \EXU/CSRControl/_0156_ ;
wire \EXU/CSRControl/_0157_ ;
wire \EXU/CSRControl/_0158_ ;
wire \EXU/CSRControl/_0159_ ;
wire \EXU/CSRControl/_0160_ ;
wire \EXU/CSRControl/_0161_ ;
wire \EXU/CSRControl/_0162_ ;
wire \EXU/CSRControl/_0163_ ;
wire \EXU/CSRControl/_0164_ ;
wire \EXU/CSRControl/_0165_ ;
wire \EXU/CSRControl/_0166_ ;
wire \EXU/CSRControl/_0167_ ;
wire \EXU/CSRControl/_0168_ ;
wire \EXU/CSRControl/_0169_ ;
wire \EXU/CSRControl/_0170_ ;
wire \EXU/CSRControl/_0171_ ;
wire \EXU/CSRControl/_0172_ ;
wire \EXU/CSRControl/_0173_ ;
wire \EXU/CSRControl/_0174_ ;
wire \EXU/CSRControl/_0175_ ;
wire \EXU/CSRControl/_0176_ ;
wire \EXU/CSRControl/_0177_ ;
wire \EXU/CSRControl/_0178_ ;
wire \EXU/CSRControl/_0179_ ;
wire \EXU/CSRControl/_0180_ ;
wire \EXU/CSRControl/_0181_ ;
wire \EXU/CSRControl/_0182_ ;
wire \EXU/CSRControl/_0183_ ;
wire \EXU/CSRControl/_0184_ ;
wire \EXU/CSRControl/_0185_ ;
wire \EXU/CSRControl/_0186_ ;
wire \EXU/CSRControl/_0187_ ;
wire \EXU/CSRControl/_0188_ ;
wire \EXU/CSRControl/_0189_ ;
wire \EXU/CSRControl/_0190_ ;
wire \EXU/CSRControl/_0191_ ;
wire \EXU/CSRControl/_0192_ ;
wire \EXU/CSRControl/_0193_ ;
wire \EXU/CSRControl/_0194_ ;
wire \EXU/CSRControl/_0195_ ;
wire \EXU/CSRControl/_0196_ ;
wire \EXU/CSRControl/_0197_ ;
wire \EXU/CSRControl/_0198_ ;
wire \EXU/CSRControl/_0199_ ;
wire \EXU/CSRControl/_0200_ ;
wire \EXU/CSRControl/_0201_ ;
wire \EXU/CSRControl/_0202_ ;
wire \EXU/CSRControl/_0203_ ;
wire \EXU/CSRControl/_0204_ ;
wire \EXU/CSRControl/_0205_ ;
wire \EXU/CSRControl/_0206_ ;
wire \EXU/CSRControl/_0207_ ;
wire \EXU/CSRControl/_0208_ ;
wire \EXU/CSRControl/_0209_ ;
wire \EXU/CSRControl/_0210_ ;
wire \EXU/CSRControl/_0211_ ;
wire \EXU/CSRControl/_0212_ ;
wire \EXU/CSRControl/_0213_ ;
wire \EXU/CSRControl/_0214_ ;
wire \EXU/CSRControl/_0215_ ;
wire \EXU/CSRControl/_0216_ ;
wire \EXU/CSRControl/_0217_ ;
wire \EXU/CSRControl/_0218_ ;
wire \EXU/CSRControl/_0219_ ;
wire \EXU/CSRControl/_0220_ ;
wire \EXU/CSRControl/_0221_ ;
wire \EXU/CSRControl/_0222_ ;
wire \EXU/CSRControl/_0223_ ;
wire \EXU/CSRControl/_0224_ ;
wire \EXU/CSRControl/_0225_ ;
wire \EXU/CSRControl/_0226_ ;
wire \EXU/CSRControl/_0227_ ;
wire \EXU/CSRControl/_0228_ ;
wire \EXU/CSRControl/_0229_ ;
wire \EXU/CSRControl/_0230_ ;
wire \EXU/CSRControl/_0231_ ;
wire \EXU/CSRControl/_0232_ ;
wire \EXU/CSRControl/_0233_ ;
wire \EXU/CSRControl/_0234_ ;
wire \EXU/CSRControl/_0235_ ;
wire \EXU/CSRControl/_0236_ ;
wire \EXU/CSRControl/_0237_ ;
wire \EXU/CSRControl/_0238_ ;
wire \EXU/CSRControl/_0239_ ;
wire \EXU/CSRControl/_0240_ ;
wire \EXU/CSRControl/_0241_ ;
wire \EXU/CSRControl/_0242_ ;
wire \EXU/CSRControl/_0243_ ;
wire \EXU/CSRControl/_0244_ ;
wire \EXU/CSRControl/_0245_ ;
wire \EXU/CSRControl/_0246_ ;
wire \EXU/CSRControl/_0247_ ;
wire \EXU/CSRControl/_0248_ ;
wire \EXU/CSRControl/_0249_ ;
wire \EXU/CSRControl/_0250_ ;
wire \EXU/CSRControl/_0251_ ;
wire \EXU/CSRControl/_0252_ ;
wire \EXU/CSRControl/_0253_ ;
wire \EXU/CSRControl/_0254_ ;
wire \EXU/CSRControl/_0255_ ;
wire \EXU/CSRControl/_0256_ ;
wire \EXU/CSRControl/_0257_ ;
wire \EXU/CSRControl/_0258_ ;
wire \EXU/CSRControl/_0259_ ;
wire \EXU/CSRControl/_0260_ ;
wire \EXU/CSRControl/_0261_ ;
wire \EXU/CSRControl/_0262_ ;
wire \EXU/CSRControl/_0263_ ;
wire \EXU/CSRControl/_0264_ ;
wire \EXU/CSRControl/_0265_ ;
wire \EXU/CSRControl/_0266_ ;
wire \EXU/CSRControl/_0267_ ;
wire \EXU/CSRControl/_0268_ ;
wire \EXU/CSRControl/_0269_ ;
wire \EXU/CSRControl/_0270_ ;
wire \EXU/CSRControl/_0271_ ;
wire \EXU/CSRControl/_0272_ ;
wire \EXU/CSRControl/_0273_ ;
wire \EXU/CSRControl/_0274_ ;
wire \EXU/CSRControl/_0275_ ;
wire \EXU/CSRControl/_0276_ ;
wire \EXU/CSRControl/_0277_ ;
wire \EXU/CSRControl/_0278_ ;
wire \EXU/CSRControl/_0279_ ;
wire \EXU/CSRControl/_0280_ ;
wire \EXU/CSRControl/_0281_ ;
wire \EXU/CSRControl/_0282_ ;
wire \EXU/CSRControl/_0283_ ;
wire \EXU/CSRControl/_0284_ ;
wire \EXU/CSRControl/_0285_ ;
wire \EXU/CSRControl/_0286_ ;
wire \EXU/CSRControl/_0287_ ;
wire \EXU/CSRControl/_0288_ ;
wire \EXU/CSRControl/_0289_ ;
wire \EXU/CSRControl/_0290_ ;
wire \EXU/CSRControl/_0291_ ;
wire \EXU/CSRControl/_0292_ ;
wire \EXU/CSRControl/_0293_ ;
wire \EXU/CSRControl/_0294_ ;
wire \EXU/CSRControl/_0295_ ;
wire \EXU/CSRControl/_0296_ ;
wire \EXU/CSRControl/_0297_ ;
wire \EXU/CSRControl/_0298_ ;
wire \EXU/CSRControl/_0299_ ;
wire \EXU/CSRControl/_0300_ ;
wire \EXU/CSRControl/_0301_ ;
wire \EXU/CSRControl/_0302_ ;
wire \EXU/CSRControl/_0303_ ;
wire \EXU/CSRControl/_0304_ ;
wire \EXU/CSRControl/_0305_ ;
wire \EXU/CSRControl/_0306_ ;
wire \EXU/CSRControl/_0307_ ;
wire \EXU/CSRControl/_0308_ ;
wire \EXU/CSRControl/_0309_ ;
wire \EXU/CSRControl/_0310_ ;
wire \EXU/CSRControl/_0311_ ;
wire \EXU/CSRControl/_0312_ ;
wire \EXU/CSRControl/_0313_ ;
wire \EXU/CSRControl/_0314_ ;
wire \EXU/CSRControl/_0315_ ;
wire \EXU/CSRControl/_0316_ ;
wire \EXU/CSRControl/_0317_ ;
wire \EXU/CSRControl/_0318_ ;
wire \EXU/CSRControl/_0319_ ;
wire \EXU/CSRControl/_0320_ ;
wire \EXU/CSRControl/_0321_ ;
wire \EXU/CSRControl/_0322_ ;
wire \EXU/CSRControl/_0323_ ;
wire \EXU/CSRControl/_0324_ ;
wire \EXU/CSRControl/_0325_ ;
wire \EXU/CSRControl/_0326_ ;
wire \EXU/CSRControl/_0327_ ;
wire \EXU/CSRControl/_0328_ ;
wire \EXU/CSRControl/_0329_ ;
wire \EXU/CSRControl/_0330_ ;
wire \EXU/CSRControl/_0331_ ;
wire \EXU/CSRControl/_0332_ ;
wire \EXU/CSRControl/_0333_ ;
wire \EXU/CSRControl/_0334_ ;
wire \EXU/CSRControl/_0335_ ;
wire \EXU/CSRControl/_0336_ ;
wire \EXU/CSRControl/_0337_ ;
wire \EXU/CSRControl/_0338_ ;
wire \EXU/CSRControl/_0339_ ;
wire \EXU/CSRControl/_0340_ ;
wire \EXU/CSRControl/_0341_ ;
wire \EXU/CSRControl/_0342_ ;
wire \EXU/CSRControl/_0343_ ;
wire \EXU/CSRControl/_0344_ ;
wire \EXU/CSRControl/_0345_ ;
wire \EXU/CSRControl/_0346_ ;
wire \EXU/CSRControl/_0347_ ;
wire \EXU/CSRControl/_0348_ ;
wire \EXU/CSRControl/_0349_ ;
wire \EXU/CSRControl/_0350_ ;
wire \EXU/CSRControl/_0351_ ;
wire \EXU/CSRControl/_0352_ ;
wire \EXU/CSRControl/_0353_ ;
wire \EXU/CSRControl/_0354_ ;
wire \EXU/CSRControl/_0355_ ;
wire \EXU/CSRControl/_0356_ ;
wire \EXU/CSRControl/_0357_ ;
wire \EXU/CSRControl/_0358_ ;
wire \EXU/CSRControl/_0359_ ;
wire \EXU/CSRControl/_0360_ ;
wire \EXU/CSRControl/_0361_ ;
wire \EXU/CSRControl/_0362_ ;
wire \EXU/CSRControl/_0363_ ;
wire \EXU/CSRControl/_0364_ ;
wire \EXU/CSRControl/_0365_ ;
wire \EXU/CSRControl/_0366_ ;
wire \EXU/CSRControl/_0367_ ;
wire \EXU/CSRControl/_0368_ ;
wire \EXU/CSRControl/_0369_ ;
wire \EXU/CSRControl/_0370_ ;
wire \EXU/CSRControl/_0371_ ;
wire \EXU/CSRControl/_0372_ ;
wire \EXU/CSRControl/_0373_ ;
wire \EXU/CSRControl/_0374_ ;
wire \EXU/CSRControl/_0375_ ;
wire \EXU/CSRControl/_0376_ ;
wire \EXU/CSRControl/_0377_ ;
wire \EXU/CSRControl/_0378_ ;
wire \EXU/CSRControl/_0379_ ;
wire \EXU/CSRControl/_0380_ ;
wire \EXU/CSRControl/_0381_ ;
wire \EXU/CSRControl/_0382_ ;
wire \EXU/CSRControl/_0383_ ;
wire \EXU/CSRControl/_0384_ ;
wire \EXU/CSRControl/_0385_ ;
wire \EXU/CSRControl/_0386_ ;
wire \EXU/CSRControl/_0387_ ;
wire \EXU/CSRControl/_0388_ ;
wire \EXU/CSRControl/_0389_ ;
wire \EXU/CSRControl/_0390_ ;
wire \EXU/CSRControl/_0391_ ;
wire \EXU/CSRControl/_0392_ ;
wire \EXU/CSRControl/_0393_ ;
wire \EXU/CSRControl/_0394_ ;
wire \EXU/CSRControl/_0395_ ;
wire \EXU/CSRControl/_0396_ ;
wire \EXU/CSRControl/_0397_ ;
wire \EXU/CSRControl/_0398_ ;
wire \EXU/CSRControl/_0399_ ;
wire \EXU/CSRControl/_0400_ ;
wire \EXU/CSRControl/_0401_ ;
wire \EXU/CSRControl/_0402_ ;
wire \EXU/CSRControl/_0403_ ;
wire \EXU/CSRControl/_0404_ ;
wire \EXU/CSRControl/_0405_ ;
wire \EXU/CSRControl/_0406_ ;
wire \EXU/CSRControl/_0407_ ;
wire \EXU/CSRControl/_0408_ ;
wire \EXU/CSRControl/_0409_ ;
wire \EXU/CSRControl/_0410_ ;
wire \EXU/CSRControl/_0411_ ;
wire \EXU/CSRControl/_0412_ ;
wire \EXU/CSRControl/_0413_ ;
wire \EXU/CSRControl/_0414_ ;
wire \EXU/CSRControl/_0415_ ;
wire \EXU/CSRControl/_0416_ ;
wire \EXU/CSRControl/_0417_ ;
wire \EXU/CSRControl/_0418_ ;
wire \EXU/CSRControl/_0419_ ;
wire \EXU/CSRControl/_0420_ ;
wire \EXU/CSRControl/_0421_ ;
wire \EXU/CSRControl/_0422_ ;
wire \EXU/CSRControl/_0423_ ;
wire \EXU/CSRControl/_0424_ ;
wire \EXU/CSRControl/_0425_ ;
wire \EXU/CSRControl/_0426_ ;
wire \EXU/CSRControl/_0427_ ;
wire \EXU/CSRControl/_0428_ ;
wire \EXU/CSRControl/_0429_ ;
wire \EXU/CSRControl/_0430_ ;
wire \EXU/CSRControl/_0431_ ;
wire \EXU/CSRControl/_0432_ ;
wire \EXU/CSRControl/_0433_ ;
wire \EXU/CSRControl/_0434_ ;
wire \EXU/CSRControl/_0435_ ;
wire \EXU/CSRControl/_0436_ ;
wire \EXU/CSRControl/_0437_ ;
wire \EXU/CSRControl/_0438_ ;
wire \EXU/CSRControl/_0439_ ;
wire \EXU/CSRControl/_0440_ ;
wire \EXU/CSRControl/_0441_ ;
wire \EXU/CSRControl/_0442_ ;
wire \EXU/CSRControl/_0443_ ;
wire \EXU/CSRControl/_0444_ ;
wire \EXU/CSRControl/_0445_ ;
wire \EXU/CSRControl/_0446_ ;
wire \EXU/CSRControl/_0447_ ;
wire \EXU/CSRControl/_0448_ ;
wire \EXU/CSRControl/_0449_ ;
wire \EXU/CSRControl/_0450_ ;
wire \EXU/CSRControl/_0451_ ;
wire \EXU/CSRControl/_0452_ ;
wire \EXU/CSRControl/_0453_ ;
wire \EXU/CSRControl/_0454_ ;
wire \EXU/CSRControl/_0455_ ;
wire \EXU/CSRControl/_0456_ ;
wire \EXU/CSRControl/_0457_ ;
wire \EXU/CSRControl/_0458_ ;
wire \EXU/CSRControl/_0459_ ;
wire \EXU/CSRControl/_0460_ ;
wire \EXU/CSRControl/_0461_ ;
wire \EXU/CSRControl/_0462_ ;
wire \EXU/CSRControl/_0463_ ;
wire \EXU/CSRControl/_0464_ ;
wire \EXU/CSRControl/_0465_ ;
wire \EXU/CSRControl/_0466_ ;
wire \EXU/CSRControl/_0467_ ;
wire \EXU/CSRControl/_0468_ ;
wire \EXU/CSRControl/_0469_ ;
wire \EXU/CSRControl/_0470_ ;
wire \EXU/CSRControl/_0471_ ;
wire \EXU/CSRControl/_0472_ ;
wire \EXU/CSRControl/_0473_ ;
wire \EXU/CSRControl/_0474_ ;
wire \EXU/CSRControl/_0475_ ;
wire \EXU/CSRControl/_0476_ ;
wire \EXU/CSRControl/_0477_ ;
wire \EXU/CSRControl/_0478_ ;
wire \EXU/CSRControl/_0479_ ;
wire \EXU/CSRControl/_0480_ ;
wire \EXU/CSRControl/_0481_ ;
wire \EXU/CSRControl/_0482_ ;
wire \EXU/CSRControl/_0483_ ;
wire \EXU/CSRControl/_0484_ ;
wire \EXU/CSRControl/_0485_ ;
wire \EXU/CSRControl/_0486_ ;
wire \EXU/CSRControl/_0487_ ;
wire \EXU/CSRControl/_0488_ ;
wire \EXU/CSRControl/_0489_ ;
wire \EXU/CSRControl/_0490_ ;
wire \EXU/CSRControl/_0491_ ;
wire \EXU/CSRControl/_0492_ ;
wire \EXU/CSRControl/_0493_ ;
wire \EXU/CSRControl/_0494_ ;
wire \EXU/CSRControl/_0495_ ;
wire \EXU/CSRControl/_0496_ ;
wire \EXU/CSRControl/_0497_ ;
wire \EXU/CSRControl/_0498_ ;
wire \EXU/CSRControl/_0499_ ;
wire \EXU/CSRControl/_0500_ ;
wire \EXU/CSRControl/_0501_ ;
wire \EXU/CSRControl/_0502_ ;
wire \EXU/CSRControl/_0503_ ;
wire \EXU/CSRControl/_0504_ ;
wire \EXU/CSRControl/_0505_ ;
wire \EXU/CSRControl/_0506_ ;
wire \EXU/CSRControl/_0507_ ;
wire \EXU/CSRControl/_0508_ ;
wire \EXU/CSRControl/_0509_ ;
wire \EXU/CSRControl/_0510_ ;
wire \EXU/CSRControl/_0511_ ;
wire \EXU/CSRControl/_0512_ ;
wire \EXU/CSRControl/_0513_ ;
wire \EXU/CSRControl/_0514_ ;
wire \EXU/CSRControl/_0515_ ;
wire \EXU/CSRControl/_0516_ ;
wire \EXU/CSRControl/_0517_ ;
wire \EXU/CSRControl/_0518_ ;
wire \EXU/CSRControl/_0519_ ;
wire \EXU/CSRControl/_0520_ ;
wire \EXU/CSRControl/_0521_ ;
wire \EXU/CSRControl/_0522_ ;
wire \EXU/CSRControl/_0523_ ;
wire \EXU/CSRControl/_0524_ ;
wire \EXU/CSRControl/_0525_ ;
wire \EXU/CSRControl/_0526_ ;
wire \EXU/CSRControl/_0527_ ;
wire \EXU/CSRControl/_0528_ ;
wire \EXU/CSRControl/_0529_ ;
wire \EXU/CSRControl/_0530_ ;
wire \EXU/CSRControl/_0531_ ;
wire \EXU/CSRControl/_0532_ ;
wire \EXU/CSRControl/_0533_ ;
wire \EXU/CSRControl/_0534_ ;
wire \EXU/CSRControl/_0535_ ;
wire \EXU/CSRControl/_0536_ ;
wire \EXU/CSRControl/_0537_ ;
wire \EXU/CSRControl/_0538_ ;
wire \EXU/CSRControl/_0539_ ;
wire \EXU/CSRControl/_0540_ ;
wire \EXU/CSRControl/_0541_ ;
wire \EXU/CSRControl/_0542_ ;
wire \EXU/CSRControl/_0543_ ;
wire \EXU/CSRControl/_0544_ ;
wire \EXU/CSRControl/_0545_ ;
wire \EXU/CSRControl/_0546_ ;
wire \EXU/CSRControl/_0547_ ;
wire \EXU/CSRControl/_0548_ ;
wire \EXU/CSRControl/_0549_ ;
wire \EXU/CSRControl/_0550_ ;
wire \EXU/CSRControl/_0551_ ;
wire \EXU/CSRControl/_0552_ ;
wire \EXU/CSRControl/_0553_ ;
wire \EXU/CSRControl/_0554_ ;
wire \EXU/CSRControl/_0555_ ;
wire \EXU/CSRControl/_0556_ ;
wire \EXU/CSRControl/_0557_ ;
wire \EXU/CSRControl/_0558_ ;
wire \EXU/CSRControl/_0559_ ;
wire \EXU/CSRControl/_0560_ ;
wire \EXU/CSRControl/_0561_ ;
wire \EXU/CSRControl/_0562_ ;
wire \EXU/CSRControl/_0563_ ;
wire \EXU/CSRControl/_0564_ ;
wire \EXU/CSRControl/_0565_ ;
wire \EXU/CSRControl/_0566_ ;
wire \EXU/CSRControl/_0567_ ;
wire \EXU/CSRControl/_0568_ ;
wire \EXU/CSRControl/_0569_ ;
wire \EXU/CSRControl/_0570_ ;
wire \EXU/CSRControl/_0571_ ;
wire \EXU/CSRControl/_0572_ ;
wire \EXU/CSRControl/_0573_ ;
wire \EXU/CSRControl/_0574_ ;
wire \EXU/CSRControl/_0575_ ;
wire \EXU/CSRControl/_0576_ ;
wire \EXU/CSRControl/_0577_ ;
wire \EXU/CSRControl/_0578_ ;
wire \EXU/CSRControl/_0579_ ;
wire \EXU/CSRControl/_0580_ ;
wire \EXU/CSRControl/_0581_ ;
wire \EXU/CSRControl/_0582_ ;
wire \EXU/CSRControl/_0583_ ;
wire \EXU/CSRControl/_0584_ ;
wire \EXU/CSRControl/_0585_ ;
wire \EXU/CSRControl/_0586_ ;
wire \EXU/CSRControl/_0587_ ;
wire \EXU/CSRControl/_0588_ ;
wire \EXU/CSRControl/_0589_ ;
wire \EXU/CSRControl/_0590_ ;
wire \EXU/CSRControl/_0591_ ;
wire \EXU/CSRControl/_0592_ ;
wire \EXU/CSRControl/_0593_ ;
wire \EXU/CSRControl/_0594_ ;
wire \EXU/CSRControl/_0595_ ;
wire \EXU/CSRControl/_0596_ ;
wire \EXU/CSRControl/_0597_ ;
wire \EXU/CSRControl/_0598_ ;
wire \EXU/CSRControl/_0599_ ;
wire \EXU/CSRControl/_0600_ ;
wire \EXU/CSRControl/_0601_ ;
wire \EXU/CSRControl/_0602_ ;
wire \EXU/CSRControl/_0603_ ;
wire \EXU/CSRControl/_0604_ ;
wire \EXU/CSRControl/_0605_ ;
wire \EXU/CSRControl/_0606_ ;
wire \EXU/CSRControl/_0607_ ;
wire \EXU/CSRControl/_0608_ ;
wire \EXU/CSRControl/_0609_ ;
wire \EXU/CSRControl/_0610_ ;
wire \EXU/CSRControl/_0611_ ;
wire \EXU/CSRControl/_0612_ ;
wire \EXU/CSRControl/_0613_ ;
wire \EXU/CSRControl/_0614_ ;
wire \EXU/CSRControl/_0615_ ;
wire \EXU/CSRControl/_0616_ ;
wire \EXU/CSRControl/_0617_ ;
wire \EXU/CSRControl/_0618_ ;
wire \EXU/CSRControl/_0619_ ;
wire \EXU/CSRControl/_0620_ ;
wire \EXU/CSRControl/_0621_ ;
wire \EXU/CSRControl/_0622_ ;
wire \EXU/CSRControl/_0623_ ;
wire \EXU/CSRControl/_0624_ ;
wire \EXU/CSRControl/_0625_ ;
wire \EXU/CSRControl/_0626_ ;
wire \EXU/CSRControl/_0627_ ;
wire \EXU/CSRControl/_0628_ ;
wire \EXU/CSRControl/_0629_ ;
wire \EXU/CSRControl/_0630_ ;
wire \EXU/CSRControl/_0631_ ;
wire \EXU/CSRControl/_0632_ ;
wire \EXU/CSRControl/_0633_ ;
wire \EXU/CSRControl/_0634_ ;
wire \EXU/CSRControl/_0635_ ;
wire \EXU/CSRControl/_0636_ ;
wire \EXU/CSRControl/_0637_ ;
wire \EXU/CSRControl/_0638_ ;
wire \EXU/CSRControl/_0639_ ;
wire \EXU/CSRControl/_0640_ ;
wire \EXU/CSRControl/_0641_ ;
wire \EXU/CSRControl/_0642_ ;
wire \EXU/CSRControl/_0643_ ;
wire \EXU/CSRControl/_0644_ ;
wire \EXU/CSRControl/_0645_ ;
wire \EXU/CSRControl/_0646_ ;
wire \EXU/CSRControl/_0647_ ;
wire \EXU/CSRControl/_0648_ ;
wire \EXU/CSRControl/_0649_ ;
wire \EXU/CSRControl/_0650_ ;
wire \EXU/CSRControl/_0651_ ;
wire \EXU/CSRControl/_0652_ ;
wire \EXU/CSRControl/_0653_ ;
wire \EXU/CSRControl/_0654_ ;
wire \EXU/CSRControl/_0655_ ;
wire \EXU/CSRControl/_0656_ ;
wire \EXU/CSRControl/_0657_ ;
wire \EXU/CSRControl/_0658_ ;
wire \EXU/CSRControl/_0659_ ;
wire \EXU/CSRControl/_0660_ ;
wire \EXU/CSRControl/_0661_ ;
wire \EXU/CSRControl/_0662_ ;
wire \EXU/CSRControl/_0663_ ;
wire \EXU/CSRControl/_0664_ ;
wire \EXU/CSRControl/_0665_ ;
wire \EXU/CSRControl/_0666_ ;
wire \EXU/CSRControl/_0667_ ;
wire \EXU/CSRControl/_0668_ ;
wire \EXU/CSRControl/_0669_ ;
wire \EXU/CSRControl/_0670_ ;
wire \EXU/CSRControl/_0671_ ;
wire \EXU/CSRControl/_0672_ ;
wire \EXU/CSRControl/_0673_ ;
wire \EXU/CSRControl/_0674_ ;
wire \EXU/CSRControl/_0675_ ;
wire \EXU/CSRControl/_0676_ ;
wire \EXU/CSRControl/_0677_ ;
wire \EXU/CSRControl/_0678_ ;
wire \EXU/CSRControl/_0679_ ;
wire \EXU/CSRControl/_0680_ ;
wire \EXU/CSRControl/_0681_ ;
wire \EXU/CSRControl/_0682_ ;
wire \EXU/CSRControl/_0683_ ;
wire \EXU/CSRControl/_0684_ ;
wire \EXU/CSRControl/_0685_ ;
wire \EXU/CSRControl/_0686_ ;
wire \EXU/CSRControl/_0687_ ;
wire \EXU/CSRControl/_0688_ ;
wire \EXU/CSRControl/_0689_ ;
wire \EXU/CSRControl/_0690_ ;
wire \EXU/CSRControl/_0691_ ;
wire \EXU/CSRControl/_0692_ ;
wire \EXU/CSRControl/_0693_ ;
wire \EXU/CSRControl/_0694_ ;
wire \EXU/CSRControl/_0695_ ;
wire \EXU/CSRControl/_0696_ ;
wire \EXU/CSRControl/_0697_ ;
wire \EXU/CSRControl/_0698_ ;
wire \EXU/CSRControl/_0699_ ;
wire \EXU/CSRControl/_0700_ ;
wire \EXU/CSRControl/_0701_ ;
wire \EXU/CSRControl/_0702_ ;
wire \EXU/CSRControl/_0703_ ;
wire \EXU/CSRControl/_0704_ ;
wire \EXU/CSRControl/_0705_ ;
wire \EXU/CSRControl/_0706_ ;
wire \EXU/CSRControl/_0707_ ;
wire \EXU/CSRControl/_0708_ ;
wire \EXU/CSRControl/_0709_ ;
wire \EXU/CSRControl/_0710_ ;
wire \EXU/CSRControl/_0711_ ;
wire \EXU/CSRControl/_0712_ ;
wire \EXU/CSRControl/_0713_ ;
wire \EXU/CSRControl/_0714_ ;
wire \EXU/CSRControl/_0715_ ;
wire \EXU/CSRControl/_0716_ ;
wire \EXU/CSRControl/_0717_ ;
wire \EXU/CSRControl/_0718_ ;
wire \EXU/CSRControl/_0719_ ;
wire \EXU/CSRControl/_0720_ ;
wire \EXU/CSRControl/_0721_ ;
wire \EXU/CSRControl/_0722_ ;
wire \EXU/CSRControl/_0723_ ;
wire \EXU/CSRControl/_0724_ ;
wire \EXU/CSRControl/_0725_ ;
wire \EXU/CSRControl/_0726_ ;
wire \EXU/CSRControl/_0727_ ;
wire \EXU/CSRControl/_0728_ ;
wire \EXU/CSRControl/_0729_ ;
wire \EXU/CSRControl/_0730_ ;
wire \EXU/CSRControl/_0731_ ;
wire \EXU/CSRControl/_0732_ ;
wire \EXU/CSRControl/_0733_ ;
wire \EXU/CSRControl/_0734_ ;
wire \EXU/CSRControl/_0735_ ;
wire \EXU/CSRControl/_0736_ ;
wire \EXU/CSRControl/_0737_ ;
wire \EXU/CSRControl/_0738_ ;
wire \EXU/CSRControl/_0739_ ;
wire \EXU/CSRControl/_0740_ ;
wire \EXU/CSRControl/_0741_ ;
wire \EXU/CSRControl/_0742_ ;
wire \EXU/CSRControl/_0743_ ;
wire \EXU/CSRControl/_0744_ ;
wire \EXU/CSRControl/_0745_ ;
wire \EXU/CSRControl/_0746_ ;
wire \EXU/CSRControl/_0747_ ;
wire \EXU/CSRControl/_0748_ ;
wire \EXU/CSRControl/_0749_ ;
wire \EXU/CSRControl/_0750_ ;
wire \EXU/CSRControl/_0751_ ;
wire \EXU/CSRControl/_0752_ ;
wire \EXU/CSRControl/_0753_ ;
wire \EXU/CSRControl/_0754_ ;
wire \EXU/CSRControl/_0755_ ;
wire \EXU/CSRControl/_0756_ ;
wire \EXU/CSRControl/_0757_ ;
wire \EXU/CSRControl/_0758_ ;
wire \EXU/CSRControl/_0759_ ;
wire \EXU/CSRControl/_0760_ ;
wire \EXU/CSRControl/_0761_ ;
wire \EXU/CSRControl/_0762_ ;
wire \EXU/CSRControl/_0763_ ;
wire \EXU/CSRControl/_0764_ ;
wire \EXU/CSRControl/_0765_ ;
wire \EXU/CSRControl/_0766_ ;
wire \EXU/CSRControl/_0767_ ;
wire \EXU/CSRControl/_0768_ ;
wire \EXU/CSRControl/_0769_ ;
wire \EXU/CSRControl/_0770_ ;
wire \EXU/CSRControl/_0771_ ;
wire \EXU/CSRControl/_0772_ ;
wire \EXU/CSRControl/_0773_ ;
wire \EXU/CSRControl/_0774_ ;
wire \EXU/CSRControl/_0775_ ;
wire \EXU/CSRControl/_0776_ ;
wire \EXU/CSRControl/_0777_ ;
wire \EXU/CSRControl/_0778_ ;
wire \EXU/CSRControl/_0779_ ;
wire \EXU/CSRControl/_0780_ ;
wire \EXU/CSRControl/_0781_ ;
wire \EXU/CSRControl/_0782_ ;
wire \EXU/CSRControl/_0783_ ;
wire \EXU/CSRControl/_0784_ ;
wire \EXU/CSRControl/_0785_ ;
wire \EXU/CSRControl/_0786_ ;
wire \EXU/CSRControl/_0787_ ;
wire \EXU/CSRControl/_0788_ ;
wire \EXU/CSRControl/_0789_ ;
wire \EXU/CSRControl/_0790_ ;
wire \EXU/CSRControl/_0791_ ;
wire \EXU/CSRControl/_0792_ ;
wire \EXU/CSRControl/_0793_ ;
wire \EXU/CSRControl/_0794_ ;
wire \EXU/CSRControl/_0795_ ;
wire \EXU/CSRControl/_0796_ ;
wire \EXU/CSRControl/_0797_ ;
wire \EXU/CSRControl/_0798_ ;
wire \EXU/CSRControl/_0799_ ;
wire \EXU/CSRControl/_0800_ ;
wire \EXU/CSRControl/_0801_ ;
wire \EXU/CSRControl/_0802_ ;
wire \EXU/CSRControl/_0803_ ;
wire \EXU/CSRControl/_0804_ ;
wire \EXU/CSRControl/_0805_ ;
wire \EXU/CSRControl/_0806_ ;
wire \EXU/CSRControl/_0807_ ;
wire \EXU/CSRControl/_0808_ ;
wire \EXU/CSRControl/_0809_ ;
wire \EXU/CSRControl/_0810_ ;
wire \EXU/CSRControl/_0811_ ;
wire \EXU/CSRControl/_0812_ ;
wire \EXU/CSRControl/_0813_ ;
wire \EXU/CSRControl/_0814_ ;
wire \EXU/CSRControl/_0815_ ;
wire \EXU/CSRControl/_0816_ ;
wire \EXU/CSRControl/_0817_ ;
wire \EXU/CSRControl/_0818_ ;
wire \EXU/CSRControl/_0819_ ;
wire \EXU/CSRControl/_0820_ ;
wire \EXU/CSRControl/_0821_ ;
wire \EXU/CSRControl/_0822_ ;
wire \EXU/CSRControl/_0823_ ;
wire \EXU/CSRControl/_0824_ ;
wire \EXU/CSRControl/_0825_ ;
wire \EXU/CSRControl/_0826_ ;
wire \EXU/CSRControl/_0827_ ;
wire \EXU/CSRControl/_0828_ ;
wire \EXU/CSRControl/_0829_ ;
wire \EXU/CSRControl/_0830_ ;
wire \EXU/CSRControl/_0831_ ;
wire \EXU/CSRControl/_0832_ ;
wire \EXU/CSRControl/_0833_ ;
wire \EXU/CSRControl/_0834_ ;
wire \EXU/CSRControl/_0835_ ;
wire \EXU/CSRControl/_0836_ ;
wire \EXU/CSRControl/_0837_ ;
wire \EXU/CSRControl/_0838_ ;
wire \EXU/CSRControl/_0839_ ;
wire \EXU/CSRControl/_0840_ ;
wire \EXU/CSRControl/_0841_ ;
wire \EXU/CSRControl/_0842_ ;
wire \EXU/CSRControl/_0843_ ;
wire \EXU/CSRControl/_0844_ ;
wire \EXU/CSRControl/_0845_ ;
wire \EXU/CSRControl/_0846_ ;
wire \EXU/CSRControl/_0847_ ;
wire \EXU/CSRControl/_0848_ ;
wire \EXU/CSRControl/_0849_ ;
wire \EXU/CSRControl/_0850_ ;
wire \EXU/CSRControl/_0851_ ;
wire \EXU/CSRControl/_0852_ ;
wire \EXU/CSRControl/_0853_ ;
wire \EXU/CSRControl/_0854_ ;
wire \EXU/CSRControl/_0855_ ;
wire \EXU/CSRControl/_0856_ ;
wire \EXU/CSRControl/_0857_ ;
wire \EXU/CSRControl/_0858_ ;
wire \EXU/CSRControl/_0859_ ;
wire \EXU/CSRControl/_0860_ ;
wire \EXU/CSRControl/_0861_ ;
wire \EXU/CSRControl/_0862_ ;
wire \EXU/CSRControl/_0863_ ;
wire \EXU/CSRControl/_0864_ ;
wire \EXU/CSRControl/_0865_ ;
wire \EXU/CSRControl/_0866_ ;
wire \EXU/CSRControl/_0867_ ;
wire \EXU/CSRControl/_0868_ ;
wire \EXU/CSRControl/_0869_ ;
wire \EXU/CSRControl/_0870_ ;
wire \EXU/CSRControl/_0871_ ;
wire \EXU/CSRControl/_0872_ ;
wire \EXU/CSRControl/_0873_ ;
wire \EXU/CSRControl/_0874_ ;
wire \EXU/CSRControl/_0875_ ;
wire \EXU/CSRControl/_0876_ ;
wire \EXU/CSRControl/_0877_ ;
wire \EXU/CSRControl/_0878_ ;
wire \EXU/CSRControl/_0879_ ;
wire \EXU/CSRControl/_0880_ ;
wire \EXU/CSRControl/_0881_ ;
wire \EXU/CSRControl/_0882_ ;
wire \EXU/CSRControl/_0883_ ;
wire \EXU/CSRControl/_0884_ ;
wire \EXU/CSRControl/_0885_ ;
wire \EXU/CSRControl/_0886_ ;
wire \EXU/CSRControl/_0887_ ;
wire \EXU/CSRControl/_0888_ ;
wire \EXU/CSRControl/_0889_ ;
wire \EXU/CSRControl/_0890_ ;
wire \EXU/CSRControl/_0891_ ;
wire \EXU/CSRControl/_0892_ ;
wire \EXU/CSRControl/_0893_ ;
wire \EXU/CSRControl/_0894_ ;
wire \EXU/CSRControl/_0895_ ;
wire \EXU/CSRControl/_0896_ ;
wire \EXU/CSRControl/_0897_ ;
wire \EXU/CSRControl/_0898_ ;
wire \EXU/CSRControl/_0899_ ;
wire \EXU/CSRControl/_0900_ ;
wire \EXU/CSRControl/_0901_ ;
wire \EXU/CSRControl/_0902_ ;
wire \EXU/CSRControl/_0903_ ;
wire \EXU/CSRControl/_0904_ ;
wire \EXU/CSRControl/_0905_ ;
wire \EXU/CSRControl/_0906_ ;
wire \EXU/CSRControl/_0907_ ;
wire \EXU/CSRControl/_0908_ ;
wire \EXU/CSRControl/_0909_ ;
wire \EXU/CSRControl/_0910_ ;
wire \EXU/CSRControl/_0911_ ;
wire \EXU/CSRControl/_0912_ ;
wire \EXU/CSRControl/_0913_ ;
wire \EXU/CSRControl/_0914_ ;
wire \EXU/CSRControl/_0915_ ;
wire \EXU/CSRControl/_0916_ ;
wire \EXU/CSRControl/_0917_ ;
wire \EXU/CSRControl/_0918_ ;
wire \EXU/CSRControl/_0919_ ;
wire \EXU/CSRControl/_0920_ ;
wire \EXU/CSRControl/_0921_ ;
wire \EXU/CSRControl/_0922_ ;
wire \EXU/CSRControl/_0923_ ;
wire \EXU/CSRControl/_0924_ ;
wire \EXU/CSRControl/_0925_ ;
wire \EXU/CSRControl/_0926_ ;
wire \EXU/CSRControl/_0927_ ;
wire \EXU/CSRControl/_0928_ ;
wire \EXU/CSRControl/_0929_ ;
wire \EXU/CSRControl/_0930_ ;
wire \EXU/CSRControl/_0931_ ;
wire \EXU/CSRControl/_0932_ ;
wire \EXU/CSRControl/_0933_ ;
wire \EXU/CSRControl/_0934_ ;
wire \EXU/CSRControl/_0935_ ;
wire \EXU/CSRControl/_0936_ ;
wire \EXU/CSRControl/_0937_ ;
wire \EXU/CSRControl/_0938_ ;
wire \EXU/CSRControl/_0939_ ;
wire \EXU/CSRControl/_0940_ ;
wire \EXU/CSRControl/_0941_ ;
wire \EXU/CSRControl/_0942_ ;
wire \EXU/CSRControl/_0943_ ;
wire \EXU/CSRControl/_0944_ ;
wire \EXU/CSRControl/_0945_ ;
wire \EXU/CSRControl/_0946_ ;
wire \EXU/CSRControl/_0947_ ;
wire \EXU/CSRControl/_0948_ ;
wire \EXU/CSRControl/_0949_ ;
wire \EXU/CSRControl/_0950_ ;
wire \EXU/CSRControl/_0951_ ;
wire \EXU/CSRControl/_0952_ ;
wire \EXU/CSRControl/_0953_ ;
wire \EXU/CSRControl/_0954_ ;
wire \EXU/CSRControl/_0955_ ;
wire \EXU/CSRControl/_0956_ ;
wire \EXU/CSRControl/_0957_ ;
wire \EXU/CSRControl/_0958_ ;
wire \EXU/CSRControl/_0959_ ;
wire \EXU/CSRControl/_0960_ ;
wire \EXU/CSRControl/_0961_ ;
wire \EXU/CSRControl/_0962_ ;
wire \EXU/CSRControl/_0963_ ;
wire \EXU/CSRControl/_0964_ ;
wire \EXU/CSRControl/_0965_ ;
wire \EXU/CSRControl/_0966_ ;
wire \EXU/CSRControl/_0967_ ;
wire \EXU/CSRControl/_0968_ ;
wire \EXU/CSRControl/_0969_ ;
wire \EXU/CSRControl/_0970_ ;
wire \EXU/CSRControl/_0971_ ;
wire \EXU/CSRControl/_0972_ ;
wire \EXU/CSRControl/_0973_ ;
wire \EXU/CSRControl/_0974_ ;
wire \EXU/CSRControl/_0975_ ;
wire \EXU/CSRControl/_0976_ ;
wire \EXU/CSRControl/_0977_ ;
wire \EXU/CSRControl/_0978_ ;
wire \EXU/CSRControl/_0979_ ;
wire \EXU/CSRControl/_0980_ ;
wire \EXU/CSRControl/_0981_ ;
wire \EXU/CSRControl/_0982_ ;
wire \EXU/CSRControl/_0983_ ;
wire \EXU/CSRControl/_0984_ ;
wire \EXU/CSRControl/_0985_ ;
wire \EXU/CSRControl/_0986_ ;
wire \EXU/CSRControl/_0987_ ;
wire \EXU/CSRControl/_0988_ ;
wire \EXU/CSRControl/_0989_ ;
wire \EXU/CSRControl/_0990_ ;
wire \EXU/CSRControl/_0991_ ;
wire \EXU/CSRControl/_0992_ ;
wire \EXU/CSRControl/_0993_ ;
wire \EXU/CSRControl/_0994_ ;
wire \EXU/CSRControl/_0995_ ;
wire \EXU/CSRControl/_0996_ ;
wire \EXU/CSRControl/_0997_ ;
wire \EXU/CSRControl/_0998_ ;
wire \EXU/CSRControl/_0999_ ;
wire \EXU/CSRControl/_1000_ ;
wire \EXU/CSRControl/_1001_ ;
wire \EXU/CSRControl/_1002_ ;
wire \EXU/CSRControl/_1003_ ;
wire \EXU/CSRControl/_1004_ ;
wire \EXU/CSRControl/_1005_ ;
wire \EXU/CSRControl/_1006_ ;
wire \EXU/CSRControl/_1007_ ;
wire \EXU/CSRControl/_1008_ ;
wire \EXU/CSRControl/_1009_ ;
wire \EXU/CSRControl/_1010_ ;
wire \EXU/CSRControl/_1011_ ;
wire \EXU/CSRControl/_1012_ ;
wire \EXU/CSRControl/_1013_ ;
wire \EXU/CSRControl/_1014_ ;
wire \EXU/CSRControl/_1015_ ;
wire \EXU/CSRControl/_1016_ ;
wire \EXU/CSRControl/_1017_ ;
wire \EXU/CSRControl/_1018_ ;
wire \EXU/CSRControl/_1019_ ;
wire \EXU/CSRControl/_1020_ ;
wire \EXU/CSRControl/_1021_ ;
wire \EXU/CSRControl/_1022_ ;
wire \EXU/CSRControl/_1023_ ;
wire \EXU/CSRControl/_1024_ ;
wire \EXU/CSRControl/_1025_ ;
wire \EXU/CSRControl/_1026_ ;
wire \EXU/CSRControl/_1027_ ;
wire \EXU/CSRControl/_1028_ ;
wire \EXU/CSRControl/_1029_ ;
wire \EXU/CSRControl/_1030_ ;
wire \EXU/CSRControl/_1031_ ;
wire \EXU/CSRControl/_1032_ ;
wire \EXU/CSRControl/_1033_ ;
wire \EXU/CSRControl/_1034_ ;
wire \EXU/CSRControl/_1035_ ;
wire \EXU/CSRControl/_1036_ ;
wire \EXU/CSRControl/_1037_ ;
wire \EXU/CSRControl/_1038_ ;
wire \EXU/CSRControl/_1039_ ;
wire \EXU/CSRControl/_1040_ ;
wire \EXU/CSRControl/_1041_ ;
wire \EXU/CSRControl/_1042_ ;
wire \EXU/CSRControl/_1043_ ;
wire \EXU/CSRControl/_1044_ ;
wire \EXU/CSRControl/_1045_ ;
wire \EXU/CSRControl/_1046_ ;
wire \EXU/CSRControl/_1047_ ;
wire \EXU/CSRControl/_1048_ ;
wire \EXU/CSRControl/_1049_ ;
wire \EXU/CSRControl/_1050_ ;
wire \EXU/CSRControl/_1051_ ;
wire \EXU/CSRControl/_1052_ ;
wire \EXU/CSRControl/_1053_ ;
wire \EXU/CSRControl/_1054_ ;
wire \EXU/CSRControl/_1055_ ;
wire \EXU/CSRControl/_1056_ ;
wire \EXU/CSRControl/_1057_ ;
wire \EXU/CSRControl/_1058_ ;
wire \EXU/CSRControl/_1059_ ;
wire \EXU/CSRControl/_1060_ ;
wire \EXU/CSRControl/_1061_ ;
wire \EXU/CSRControl/_1062_ ;
wire \EXU/CSRControl/_1063_ ;
wire \EXU/CSRControl/_1064_ ;
wire \EXU/CSRControl/_1065_ ;
wire \EXU/CSRControl/_1066_ ;
wire \EXU/CSRControl/_1067_ ;
wire \EXU/CSRControl/_1068_ ;
wire \EXU/CSRControl/_1069_ ;
wire \EXU/CSRControl/_1070_ ;
wire \EXU/CSRControl/_1071_ ;
wire \EXU/CSRControl/_1072_ ;
wire \EXU/CSRControl/_1073_ ;
wire \EXU/CSRControl/_1074_ ;
wire \EXU/CSRControl/_1075_ ;
wire \EXU/CSRControl/_1076_ ;
wire \EXU/CSRControl/_1077_ ;
wire \EXU/CSRControl/_1078_ ;
wire \EXU/CSRControl/_1079_ ;
wire \EXU/CSRControl/_1080_ ;
wire \EXU/CSRControl/_1081_ ;
wire \EXU/CSRControl/_1082_ ;
wire \EXU/CSRControl/_1083_ ;
wire \EXU/CSRControl/_1084_ ;
wire \EXU/CSRControl/_1085_ ;
wire \EXU/CSRControl/_1086_ ;
wire \EXU/CSRControl/_1087_ ;
wire \EXU/CSRControl/_1088_ ;
wire \EXU/CSRControl/_1089_ ;
wire \EXU/CSRControl/_1090_ ;
wire \EXU/CSRControl/_1091_ ;
wire \EXU/CSRControl/_1092_ ;
wire \EXU/CSRControl/_1093_ ;
wire \EXU/CSRControl/_1094_ ;
wire \EXU/CSRControl/_1095_ ;
wire \EXU/CSRControl/_1096_ ;
wire \EXU/CSRControl/_1097_ ;
wire \EXU/CSRControl/_1098_ ;
wire \EXU/CSRControl/_1099_ ;
wire \EXU/CSRControl/_1100_ ;
wire \EXU/CSRControl/_1101_ ;
wire \EXU/CSRControl/_1102_ ;
wire \EXU/CSRControl/_1103_ ;
wire \EXU/CSRControl/_1104_ ;
wire \EXU/CSRControl/_1105_ ;
wire \EXU/CSRControl/_1106_ ;
wire \EXU/CSRControl/_1107_ ;
wire \EXU/CSRControl/_1108_ ;
wire \EXU/CSRControl/_1109_ ;
wire \EXU/CSRControl/_1110_ ;
wire \EXU/CSRControl/_1111_ ;
wire \EXU/CSRControl/_1112_ ;
wire \EXU/CSRControl/_1113_ ;
wire \EXU/CSRControl/_1114_ ;
wire \EXU/CSRControl/_1115_ ;
wire \EXU/CSRControl/_1116_ ;
wire \EXU/CSRControl/_1117_ ;
wire \EXU/CSRControl/_1118_ ;
wire \EXU/CSRControl/_1119_ ;
wire \EXU/CSRControl/_1120_ ;
wire \EXU/CSRControl/_1121_ ;
wire \EXU/CSRControl/_1122_ ;
wire \EXU/CSRControl/_1123_ ;
wire \EXU/CSRControl/_1124_ ;
wire \EXU/CSRControl/_1125_ ;
wire \EXU/CSRControl/_1126_ ;
wire \EXU/CSRControl/_1127_ ;
wire \EXU/CSRControl/_1128_ ;
wire \EXU/CSRControl/_1129_ ;
wire \EXU/CSRControl/_1130_ ;
wire \EXU/CSRControl/_1131_ ;
wire \EXU/CSRControl/_1132_ ;
wire \EXU/CSRControl/_1133_ ;
wire \EXU/CSRControl/_1134_ ;
wire \EXU/CSRControl/_1135_ ;
wire \EXU/CSRControl/_1136_ ;
wire \EXU/CSRControl/_1137_ ;
wire \EXU/CSRControl/_1138_ ;
wire \EXU/CSRControl/_1139_ ;
wire \EXU/CSRControl/_1140_ ;
wire \EXU/CSRControl/_1141_ ;
wire \EXU/CSRControl/_1142_ ;
wire \EXU/CSRControl/_1143_ ;
wire \EXU/CSRControl/_1144_ ;
wire \EXU/CSRControl/_1145_ ;
wire \EXU/CSRControl/_1146_ ;
wire \EXU/CSRControl/_1147_ ;
wire \EXU/CSRControl/_1148_ ;
wire \EXU/CSRControl/_1149_ ;
wire \EXU/CSRControl/_1150_ ;
wire \EXU/CSRControl/_1151_ ;
wire \EXU/CSRControl/_1152_ ;
wire \EXU/CSRControl/_1153_ ;
wire \EXU/CSRControl/_1154_ ;
wire \EXU/CSRControl/_1155_ ;
wire \EXU/CSRControl/_1156_ ;
wire \EXU/CSRControl/_1157_ ;
wire \EXU/CSRControl/_1158_ ;
wire \EXU/CSRControl/_1159_ ;
wire \EXU/CSRControl/_1160_ ;
wire \EXU/CSRControl/_1161_ ;
wire \EXU/CSRControl/_1162_ ;
wire \EXU/CSRControl/_1163_ ;
wire \EXU/CSRControl/_1164_ ;
wire \EXU/CSRControl/_1165_ ;
wire \EXU/CSRControl/_1166_ ;
wire \EXU/CSRControl/_1167_ ;
wire \EXU/CSRControl/_1168_ ;
wire \EXU/CSRControl/_1169_ ;
wire \EXU/CSRControl/_1170_ ;
wire \EXU/CSRControl/_1171_ ;
wire \EXU/CSRControl/_1172_ ;
wire \EXU/CSRControl/_1173_ ;
wire \EXU/CSRControl/_1174_ ;
wire \EXU/CSRControl/_1175_ ;
wire \EXU/CSRControl/_1176_ ;
wire \EXU/CSRControl/_1177_ ;
wire \EXU/CSRControl/_1178_ ;
wire \EXU/CSRControl/_1179_ ;
wire \EXU/CSRControl/_1180_ ;
wire \EXU/CSRControl/_1181_ ;
wire \EXU/CSRControl/_1182_ ;
wire \EXU/CSRControl/_1183_ ;
wire \EXU/CSRControl/_1184_ ;
wire \EXU/CSRControl/_1185_ ;
wire \EXU/CSRControl/_1186_ ;
wire \EXU/CSRControl/_1187_ ;
wire \EXU/CSRControl/_1188_ ;
wire \EXU/CSRControl/_1189_ ;
wire \EXU/CSRControl/_1190_ ;
wire \EXU/CSRControl/_1191_ ;
wire \EXU/CSRControl/_1192_ ;
wire \EXU/CSRControl/_1193_ ;
wire \EXU/CSRControl/_1194_ ;
wire \EXU/CSRControl/_1195_ ;
wire \EXU/CSRControl/_1196_ ;
wire \EXU/CSRControl/_1197_ ;
wire \EXU/CSRControl/_1198_ ;
wire \EXU/CSRControl/_1199_ ;
wire \EXU/CSRControl/_1200_ ;
wire \EXU/CSRControl/_1201_ ;
wire \EXU/CSRControl/_1202_ ;
wire \EXU/CSRControl/_1203_ ;
wire \EXU/CSRControl/_1204_ ;
wire \EXU/CSRControl/_1205_ ;
wire \EXU/CSRControl/_1206_ ;
wire \EXU/CSRControl/_1207_ ;
wire \EXU/CSRControl/_1208_ ;
wire \EXU/CSRControl/_1209_ ;
wire \EXU/CSRControl/_1210_ ;
wire \EXU/CSRControl/_1211_ ;
wire \EXU/CSRControl/_1212_ ;
wire \EXU/CSRControl/_1213_ ;
wire \EXU/CSRControl/_1214_ ;
wire \EXU/CSRControl/_1215_ ;
wire \EXU/CSRControl/_1216_ ;
wire \EXU/CSRControl/_1217_ ;
wire \EXU/CSRControl/_1218_ ;
wire \EXU/CSRControl/_1219_ ;
wire \EXU/CSRControl/_1220_ ;
wire \EXU/CSRControl/_1221_ ;
wire \EXU/CSRControl/_1222_ ;
wire \EXU/CSRControl/_1223_ ;
wire \EXU/CSRControl/_1224_ ;
wire \EXU/CSRControl/_1225_ ;
wire \EXU/CSRControl/_1226_ ;
wire \EXU/CSRControl/_1227_ ;
wire \EXU/CSRControl/_1228_ ;
wire \EXU/CSRControl/_1229_ ;
wire \EXU/CSRControl/_1230_ ;
wire \EXU/CSRControl/_1231_ ;
wire \EXU/CSRControl/_1232_ ;
wire \EXU/CSRControl/_1233_ ;
wire \EXU/CSRControl/_1234_ ;
wire \EXU/CSRControl/_1235_ ;
wire \EXU/CSRControl/_1236_ ;
wire \EXU/CSRControl/_1237_ ;
wire \EXU/CSRControl/_1238_ ;
wire \EXU/CSRControl/_1239_ ;
wire \EXU/CSRControl/_1240_ ;
wire \EXU/CSRControl/_1241_ ;
wire \EXU/CSRControl/_1242_ ;
wire \EXU/CSRControl/_1243_ ;
wire \EXU/CSRControl/_1244_ ;
wire \EXU/CSRControl/_1245_ ;
wire \EXU/CSRControl/_1246_ ;
wire \EXU/CSRControl/_1247_ ;
wire \EXU/CSRControl/_1248_ ;
wire \EXU/CSRControl/_1249_ ;
wire \EXU/CSRControl/_1250_ ;
wire \EXU/CSRControl/_1251_ ;
wire \EXU/CSRControl/_1252_ ;
wire \EXU/CSRControl/_1253_ ;
wire \EXU/CSRControl/_1254_ ;
wire \EXU/CSRControl/_1255_ ;
wire \EXU/CSRControl/_1256_ ;
wire \EXU/CSRControl/_1257_ ;
wire \EXU/CSRControl/_1258_ ;
wire \EXU/CSRControl/_1259_ ;
wire \EXU/CSRControl/_1260_ ;
wire \EXU/CSRControl/_1261_ ;
wire \EXU/CSRControl/_1262_ ;
wire \EXU/CSRControl/_1263_ ;
wire \EXU/CSRControl/_1264_ ;
wire \EXU/CSRControl/_1265_ ;
wire \EXU/CSRControl/_1266_ ;
wire \EXU/CSRControl/_1267_ ;
wire \EXU/CSRControl/_1268_ ;
wire \EXU/CSRControl/_1269_ ;
wire \EXU/CSRControl/_1270_ ;
wire \EXU/CSRControl/_1271_ ;
wire \EXU/CSRControl/_1272_ ;
wire \EXU/CSRControl/_1273_ ;
wire \EXU/CSRControl/_1274_ ;
wire \EXU/CSRControl/_1275_ ;
wire \EXU/CSRControl/_1276_ ;
wire \EXU/CSRControl/_1277_ ;
wire \EXU/CSRControl/_1278_ ;
wire \EXU/CSRControl/_1279_ ;
wire \EXU/CSRControl/_1280_ ;
wire \EXU/CSRControl/_1281_ ;
wire \EXU/CSRControl/_1282_ ;
wire \EXU/CSRControl/_1283_ ;
wire \EXU/CSRControl/_1284_ ;
wire \EXU/CSRControl/_1285_ ;
wire \EXU/CSRControl/_1286_ ;
wire \EXU/CSRControl/_1287_ ;
wire \EXU/CSRControl/_1288_ ;
wire \EXU/CSRControl/_1289_ ;
wire \EXU/CSRControl/_1290_ ;
wire \EXU/CSRControl/_1291_ ;
wire \EXU/CSRControl/_1292_ ;
wire \EXU/CSRControl/_1293_ ;
wire \EXU/CSRControl/_1294_ ;
wire \EXU/CSRControl/_1295_ ;
wire \EXU/CSRControl/_1296_ ;
wire \EXU/CSRControl/_1297_ ;
wire \EXU/CSRControl/_1298_ ;
wire \EXU/CSRControl/_1299_ ;
wire \EXU/CSRControl/_1300_ ;
wire \EXU/CSRControl/_1301_ ;
wire \EXU/CSRControl/_1302_ ;
wire \EXU/CSRControl/_1303_ ;
wire \EXU/CSRControl/_1304_ ;
wire \EXU/CSRControl/_1305_ ;
wire \EXU/CSRControl/_1306_ ;
wire \EXU/CSRControl/_1307_ ;
wire \EXU/CSRControl/_1308_ ;
wire \EXU/CSRControl/_1309_ ;
wire \EXU/CSRControl/_1310_ ;
wire \EXU/CSRControl/_1311_ ;
wire \EXU/CSRControl/_1312_ ;
wire \EXU/CSRControl/_1313_ ;
wire \EXU/CSRControl/_1314_ ;
wire \EXU/CSRControl/_1315_ ;
wire \EXU/CSRControl/_1316_ ;
wire \EXU/CSRControl/_1317_ ;
wire \EXU/CSRControl/_1318_ ;
wire \EXU/CSRControl/_1319_ ;
wire \EXU/CSRControl/_1320_ ;
wire \EXU/CSRControl/_1321_ ;
wire \EXU/CSRControl/_1322_ ;
wire \EXU/CSRControl/_1323_ ;
wire \EXU/CSRControl/_1324_ ;
wire \EXU/CSRControl/_1325_ ;
wire \EXU/CSRControl/_1326_ ;
wire \EXU/CSRControl/_1327_ ;
wire \EXU/CSRControl/_1328_ ;
wire \EXU/CSRControl/_1329_ ;
wire \EXU/CSRControl/_1330_ ;
wire \EXU/CSRControl/_1331_ ;
wire \EXU/CSRControl/_1332_ ;
wire \EXU/CSRControl/_1333_ ;
wire \EXU/CSRControl/_1334_ ;
wire \EXU/CSRControl/_1335_ ;
wire \EXU/CSRControl/_1336_ ;
wire \EXU/CSRControl/_1337_ ;
wire \EXU/CSRControl/_1338_ ;
wire \EXU/CSRControl/_1339_ ;
wire \EXU/CSRControl/_1340_ ;
wire \EXU/CSRControl/_1341_ ;
wire \EXU/CSRControl/_1342_ ;
wire \EXU/CSRControl/_1343_ ;
wire \EXU/CSRControl/_1344_ ;
wire \EXU/CSRControl/_1345_ ;
wire \EXU/CSRControl/_1346_ ;
wire \EXU/CSRControl/_1347_ ;
wire \EXU/CSRControl/_1348_ ;
wire \EXU/CSRControl/_1349_ ;
wire \EXU/CSRControl/_1350_ ;
wire \EXU/CSRControl/_1351_ ;
wire \EXU/CSRControl/_1352_ ;
wire \EXU/CSRControl/_1353_ ;
wire \EXU/CSRControl/_1354_ ;
wire \EXU/CSRControl/_1355_ ;
wire \EXU/CSRControl/_1356_ ;
wire \EXU/CSRControl/_1357_ ;
wire \EXU/CSRControl/_1358_ ;
wire \EXU/CSRControl/_1359_ ;
wire \EXU/CSRControl/_1360_ ;
wire \EXU/CSRControl/_1361_ ;
wire \EXU/CSRControl/_1362_ ;
wire \EXU/CSRControl/_1363_ ;
wire \EXU/CSRControl/_1364_ ;
wire \EXU/CSRControl/_1365_ ;
wire \EXU/CSRControl/_1366_ ;
wire \EXU/CSRControl/_1367_ ;
wire \EXU/CSRControl/_1368_ ;
wire \EXU/CSRControl/_1369_ ;
wire \EXU/CSRControl/_1370_ ;
wire \EXU/CSRControl/_1371_ ;
wire \EXU/CSRControl/_1372_ ;
wire \EXU/CSRControl/_1373_ ;
wire \EXU/CSRControl/_1374_ ;
wire \EXU/CSRControl/_1375_ ;
wire \EXU/CSRControl/_1376_ ;
wire \EXU/CSRControl/_1377_ ;
wire \EXU/CSRControl/_1378_ ;
wire \EXU/CSRControl/_1379_ ;
wire \EXU/CSRControl/_1380_ ;
wire \EXU/CSRControl/_1381_ ;
wire \EXU/CSRControl/_1382_ ;
wire \EXU/CSRControl/_1383_ ;
wire \EXU/CSRControl/_1384_ ;
wire \EXU/CSRControl/_1385_ ;
wire \EXU/CSRControl/_1386_ ;
wire \EXU/CSRControl/_1387_ ;
wire \EXU/CSRControl/_1388_ ;
wire \EXU/CSRControl/_1389_ ;
wire \EXU/CSRControl/_1390_ ;
wire \EXU/CSRControl/_1391_ ;
wire \EXU/CSRControl/_1392_ ;
wire \EXU/CSRControl/_1393_ ;
wire \EXU/CSRControl/_1394_ ;
wire \EXU/CSRControl/_1395_ ;
wire \EXU/CSRControl/_1396_ ;
wire \EXU/CSRControl/_1397_ ;
wire \EXU/CSRControl/_1398_ ;
wire \EXU/CSRControl/_1399_ ;
wire \EXU/CSRControl/_1400_ ;
wire \EXU/CSRControl/_1401_ ;
wire \EXU/CSRControl/_1402_ ;
wire \EXU/CSRControl/_1403_ ;
wire \EXU/CSRControl/_1404_ ;
wire \EXU/CSRControl/_1405_ ;
wire \EXU/CSRControl/_1406_ ;
wire \EXU/CSRControl/_1407_ ;
wire \EXU/CSRControl/_1408_ ;
wire \EXU/CSRControl/_1409_ ;
wire \EXU/CSRControl/_1410_ ;
wire \EXU/CSRControl/_1411_ ;
wire \EXU/CSRControl/_1412_ ;
wire \EXU/CSRControl/_1413_ ;
wire \EXU/CSRControl/_1414_ ;
wire \EXU/CSRControl/_1415_ ;
wire \EXU/CSRControl/_1416_ ;
wire \EXU/CSRControl/_1417_ ;
wire \EXU/CSRControl/_1418_ ;
wire \EXU/CSRControl/_1419_ ;
wire \EXU/CSRControl/_1420_ ;
wire \EXU/CSRControl/_1421_ ;
wire \EXU/CSRControl/_1422_ ;
wire \EXU/CSRControl/_1423_ ;
wire \EXU/CSRControl/_1424_ ;
wire \EXU/CSRControl/_1425_ ;
wire \EXU/CSRControl/_1426_ ;
wire \EXU/CSRControl/_1427_ ;
wire \EXU/CSRControl/_1428_ ;
wire \EXU/CSRControl/_1429_ ;
wire \EXU/CSRControl/_1430_ ;
wire \EXU/CSRControl/_1431_ ;
wire \EXU/CSRControl/_1432_ ;
wire \EXU/CSRControl/_1433_ ;
wire \EXU/CSRControl/_1434_ ;
wire \EXU/CSRControl/_1435_ ;
wire \EXU/CSRControl/_1436_ ;
wire \EXU/CSRControl/_1437_ ;
wire \EXU/CSRControl/_1438_ ;
wire \EXU/CSRControl/_1439_ ;
wire \EXU/CSRControl/_1440_ ;
wire \EXU/CSRControl/_1441_ ;
wire \EXU/CSRControl/_1442_ ;
wire \EXU/CSRControl/_1443_ ;
wire \EXU/CSRControl/_1444_ ;
wire \EXU/CSRControl/_1445_ ;
wire \EXU/CSRControl/_1446_ ;
wire \EXU/CSRControl/_1447_ ;
wire \EXU/CSRControl/_1448_ ;
wire \EXU/CSRControl/_1449_ ;
wire \EXU/CSRControl/_1450_ ;
wire \EXU/CSRControl/_1451_ ;
wire \EXU/CSRControl/_1452_ ;
wire \EXU/CSRControl/_1453_ ;
wire \EXU/CSRControl/_1454_ ;
wire \EXU/CSRControl/_1455_ ;
wire \EXU/CSRControl/_1456_ ;
wire \EXU/CSRControl/_1457_ ;
wire \EXU/CSRControl/_1458_ ;
wire \EXU/CSRControl/_1459_ ;
wire \EXU/CSRControl/_1460_ ;
wire \EXU/CSRControl/_1461_ ;
wire \EXU/CSRControl/_1462_ ;
wire \EXU/CSRControl/_1463_ ;
wire \EXU/CSRControl/_1464_ ;
wire \EXU/CSRControl/_1465_ ;
wire \EXU/CSRControl/_1466_ ;
wire \EXU/CSRControl/_1467_ ;
wire \EXU/CSRControl/_1468_ ;
wire \EXU/CSRControl/_1469_ ;
wire \EXU/CSRControl/_1470_ ;
wire \EXU/CSRControl/_1471_ ;
wire \EXU/CSRControl/_1472_ ;
wire \EXU/CSRControl/_1473_ ;
wire \EXU/CSRControl/_1474_ ;
wire \EXU/CSRControl/_1475_ ;
wire \EXU/CSRControl/_1476_ ;
wire \EXU/CSRControl/_1477_ ;
wire \EXU/CSRControl/_1478_ ;
wire \EXU/CSRControl/_1479_ ;
wire \EXU/CSRControl/_1480_ ;
wire \EXU/CSRControl/_1481_ ;
wire \EXU/CSRControl/_1482_ ;
wire \EXU/CSRControl/_1483_ ;
wire \EXU/CSRControl/_1484_ ;
wire \EXU/CSRControl/_1485_ ;
wire \EXU/CSRControl/_1486_ ;
wire \EXU/CSRControl/_1487_ ;
wire \EXU/CSRControl/_1488_ ;
wire \EXU/CSRControl/_1489_ ;
wire \EXU/CSRControl/_1490_ ;
wire \EXU/CSRControl/_1491_ ;
wire \EXU/CSRControl/_1492_ ;
wire \EXU/CSRControl/_1493_ ;
wire \EXU/CSRControl/_1494_ ;
wire \EXU/CSRControl/_1495_ ;
wire \EXU/CSRControl/_1496_ ;
wire \EXU/CSRControl/_1497_ ;
wire \EXU/CSRControl/_1498_ ;
wire \EXU/CSRControl/_1499_ ;
wire \EXU/CSRControl/_1500_ ;
wire \EXU/CSRControl/_1501_ ;
wire \EXU/CSRControl/_1502_ ;
wire \EXU/CSRControl/_1503_ ;
wire \EXU/CSRControl/_1504_ ;
wire \EXU/CSRControl/_1505_ ;
wire \EXU/CSRControl/_1506_ ;
wire \EXU/CSRControl/_1507_ ;
wire \EXU/CSRControl/_1508_ ;
wire \EXU/CSRControl/_1509_ ;
wire \EXU/CSRControl/_1510_ ;
wire \EXU/CSRControl/_1511_ ;
wire \EXU/CSRControl/_1512_ ;
wire \EXU/CSRControl/_1513_ ;
wire \EXU/CSRControl/_1514_ ;
wire \EXU/CSRControl/_1515_ ;
wire \EXU/CSRControl/_1516_ ;
wire \EXU/CSRControl/_1517_ ;
wire \EXU/CSRControl/_1518_ ;
wire \EXU/CSRControl/_1519_ ;
wire \EXU/CSRControl/_1520_ ;
wire \EXU/CSRControl/_1521_ ;
wire \EXU/CSRControl/_1522_ ;
wire \EXU/CSRControl/_1523_ ;
wire \EXU/CSRControl/_1524_ ;
wire \EXU/CSRControl/_1525_ ;
wire \EXU/CSRControl/_1526_ ;
wire \EXU/CSRControl/_1527_ ;
wire \EXU/CSRControl/_1528_ ;
wire \EXU/CSRControl/_1529_ ;
wire \EXU/CSRControl/_1530_ ;
wire \EXU/CSRControl/_1531_ ;
wire \EXU/CSRControl/_1532_ ;
wire \EXU/CSRControl/_1533_ ;
wire \EXU/CSRControl/_1534_ ;
wire \EXU/CSRControl/_1535_ ;
wire \EXU/CSRControl/_1536_ ;
wire \EXU/CSRControl/_1537_ ;
wire \EXU/CSRControl/_1538_ ;
wire \EXU/CSRControl/_1539_ ;
wire \EXU/CSRControl/_1540_ ;
wire \EXU/CSRControl/_1541_ ;
wire \EXU/CSRControl/_1542_ ;
wire \EXU/CSRControl/_1543_ ;
wire \EXU/CSRControl/_1544_ ;
wire \EXU/CSRControl/_1545_ ;
wire \EXU/CSRControl/_1546_ ;
wire \EXU/CSRControl/_1547_ ;
wire \EXU/CSRControl/_1548_ ;
wire \EXU/CSRControl/_1549_ ;
wire \EXU/CSRControl/_1550_ ;
wire \EXU/CSRControl/_1551_ ;
wire \EXU/CSRControl/_1552_ ;
wire \EXU/CSRControl/_1553_ ;
wire \EXU/CSRControl/_1554_ ;
wire \EXU/CSRControl/_1555_ ;
wire \EXU/CSRControl/_1556_ ;
wire \EXU/CSRControl/_1557_ ;
wire \EXU/CSRControl/_1558_ ;
wire \EXU/CSRControl/_1559_ ;
wire \EXU/CSRControl/_1560_ ;
wire \EXU/CSRControl/_1561_ ;
wire \EXU/CSRControl/_1562_ ;
wire \EXU/CSRControl/_1563_ ;
wire \EXU/CSRControl/_1564_ ;
wire \EXU/CSRControl/_1565_ ;
wire \EXU/CSRControl/_1566_ ;
wire \EXU/CSRControl/_1567_ ;
wire \EXU/CSRControl/_1568_ ;
wire \EXU/CSRControl/_1569_ ;
wire \EXU/CSRControl/_1570_ ;
wire \EXU/CSRControl/_1571_ ;
wire \EXU/CSRControl/_1572_ ;
wire \EXU/CSRControl/_1573_ ;
wire \EXU/CSRControl/_1574_ ;
wire \EXU/CSRControl/_1575_ ;
wire \EXU/CSRControl/_1576_ ;
wire \EXU/CSRControl/_1577_ ;
wire \EXU/CSRControl/_1578_ ;
wire \EXU/CSRControl/_1579_ ;
wire \EXU/CSRControl/_1580_ ;
wire \EXU/CSRControl/_1581_ ;
wire \EXU/CSRControl/_1582_ ;
wire \EXU/CSRControl/_1583_ ;
wire \EXU/CSRControl/_1584_ ;
wire \EXU/CSRControl/_1585_ ;
wire \EXU/CSRControl/_1586_ ;
wire \EXU/CSRControl/_1587_ ;
wire \EXU/CSRControl/_1588_ ;
wire \EXU/CSRControl/_1589_ ;
wire \EXU/CSRControl/_1590_ ;
wire \EXU/CSRControl/_1591_ ;
wire \EXU/CSRControl/_1592_ ;
wire \EXU/CSRControl/_1593_ ;
wire \EXU/CSRControl/_1594_ ;
wire \EXU/CSRControl/_1595_ ;
wire \EXU/CSRControl/_1596_ ;
wire \EXU/CSRControl/_1597_ ;
wire \EXU/CSRControl/_1598_ ;
wire \EXU/CSRControl/_1599_ ;
wire \EXU/CSRControl/_1600_ ;
wire \EXU/CSRControl/_1601_ ;
wire \EXU/CSRControl/_1602_ ;
wire \EXU/CSRControl/_1603_ ;
wire \EXU/CSRControl/_1604_ ;
wire \EXU/CSRControl/_1605_ ;
wire \EXU/CSRControl/_1606_ ;
wire \EXU/CSRControl/_1607_ ;
wire \EXU/CSRControl/_1608_ ;
wire \EXU/CSRControl/_1609_ ;
wire \EXU/CSRControl/_1610_ ;
wire \EXU/CSRControl/_1611_ ;
wire \EXU/CSRControl/_1612_ ;
wire \EXU/CSRControl/_1613_ ;
wire \EXU/CSRControl/_1614_ ;
wire \EXU/CSRControl/_1615_ ;
wire \EXU/CSRControl/_1616_ ;
wire \EXU/CSRControl/_1617_ ;
wire \EXU/CSRControl/_1618_ ;
wire \EXU/CSRControl/_1619_ ;
wire \EXU/CSRControl/_1620_ ;
wire \EXU/CSRControl/_1621_ ;
wire \EXU/CSRControl/_1622_ ;
wire \EXU/CSRControl/_1623_ ;
wire \EXU/CSRControl/_1624_ ;
wire \EXU/CSRControl/_1625_ ;
wire \EXU/CSRControl/_1626_ ;
wire \EXU/CSRControl/_1627_ ;
wire \EXU/CSRControl/_1628_ ;
wire \EXU/CSRControl/_1629_ ;
wire \EXU/CSRControl/_1630_ ;
wire \EXU/CSRControl/_1631_ ;
wire \EXU/CSRControl/_1632_ ;
wire \EXU/CSRControl/_1633_ ;
wire \IDU/_000_ ;
wire \IDU/_001_ ;
wire \IDU/_002_ ;
wire \IDU/_003_ ;
wire \IDU/_004_ ;
wire \IDU/_005_ ;
wire \IDU/_006_ ;
wire \IDU/_007_ ;
wire \IDU/_008_ ;
wire \IDU/_009_ ;
wire \IDU/_010_ ;
wire \IDU/_Control_io_isEnd ;
wire \IDU/Control/_000_ ;
wire \IDU/Control/_001_ ;
wire \IDU/Control/_002_ ;
wire \IDU/Control/_003_ ;
wire \IDU/Control/_004_ ;
wire \IDU/Control/_005_ ;
wire \IDU/Control/_006_ ;
wire \IDU/Control/_007_ ;
wire \IDU/Control/_008_ ;
wire \IDU/Control/_009_ ;
wire \IDU/Control/_010_ ;
wire \IDU/Control/_011_ ;
wire \IDU/Control/_012_ ;
wire \IDU/Control/_013_ ;
wire \IDU/Control/_014_ ;
wire \IDU/Control/_015_ ;
wire \IDU/Control/_016_ ;
wire \IDU/Control/_017_ ;
wire \IDU/Control/_018_ ;
wire \IDU/Control/_019_ ;
wire \IDU/Control/_020_ ;
wire \IDU/Control/_021_ ;
wire \IDU/Control/_022_ ;
wire \IDU/Control/_023_ ;
wire \IDU/Control/_024_ ;
wire \IDU/Control/_025_ ;
wire \IDU/Control/_026_ ;
wire \IDU/Control/_027_ ;
wire \IDU/Control/_028_ ;
wire \IDU/Control/_029_ ;
wire \IDU/Control/_030_ ;
wire \IDU/Control/_031_ ;
wire \IDU/Control/_032_ ;
wire \IDU/Control/_033_ ;
wire \IDU/Control/_034_ ;
wire \IDU/Control/_035_ ;
wire \IDU/Control/_036_ ;
wire \IDU/Control/_037_ ;
wire \IDU/Control/_038_ ;
wire \IDU/Control/_039_ ;
wire \IDU/Control/_040_ ;
wire \IDU/Control/_041_ ;
wire \IDU/Control/_042_ ;
wire \IDU/Control/_043_ ;
wire \IDU/Control/_044_ ;
wire \IDU/Control/_045_ ;
wire \IDU/Control/_046_ ;
wire \IDU/Control/_047_ ;
wire \IDU/Control/_048_ ;
wire \IDU/Control/_049_ ;
wire \IDU/Control/_050_ ;
wire \IDU/Control/_051_ ;
wire \IDU/Control/_052_ ;
wire \IDU/Control/_053_ ;
wire \IDU/Control/_054_ ;
wire \IDU/Control/_055_ ;
wire \IDU/Control/_056_ ;
wire \IDU/Control/_057_ ;
wire \IDU/Control/_058_ ;
wire \IDU/Control/_059_ ;
wire \IDU/Control/_060_ ;
wire \IDU/Control/_061_ ;
wire \IDU/Control/_062_ ;
wire \IDU/Control/_063_ ;
wire \IDU/Control/_064_ ;
wire \IDU/Control/_065_ ;
wire \IDU/Control/_066_ ;
wire \IDU/Control/_067_ ;
wire \IDU/Control/_068_ ;
wire \IDU/Control/_069_ ;
wire \IDU/Control/_070_ ;
wire \IDU/Control/_071_ ;
wire \IDU/Control/_072_ ;
wire \IDU/Control/_073_ ;
wire \IDU/Control/_074_ ;
wire \IDU/Control/_075_ ;
wire \IDU/Control/_076_ ;
wire \IDU/Control/_077_ ;
wire \IDU/Control/_078_ ;
wire \IDU/Control/_079_ ;
wire \IDU/Control/_080_ ;
wire \IDU/Control/_081_ ;
wire \IDU/Control/_082_ ;
wire \IDU/Control/_083_ ;
wire \IDU/Control/_084_ ;
wire \IDU/Control/_085_ ;
wire \IDU/Control/_086_ ;
wire \IDU/Control/_087_ ;
wire \IDU/Control/_088_ ;
wire \IDU/Control/_089_ ;
wire \IDU/Control/_090_ ;
wire \IDU/Control/_091_ ;
wire \IDU/Control/_092_ ;
wire \IDU/Control/_093_ ;
wire \IDU/Control/_094_ ;
wire \IDU/Control/_095_ ;
wire \IDU/Control/_096_ ;
wire \IDU/Control/_097_ ;
wire \IDU/Control/_098_ ;
wire \IDU/Control/_099_ ;
wire \IDU/Control/_100_ ;
wire \IDU/Control/_101_ ;
wire \IDU/Control/_102_ ;
wire \IDU/Control/_103_ ;
wire \IDU/Control/_104_ ;
wire \IDU/Control/_105_ ;
wire \IDU/Control/_106_ ;
wire \IDU/Control/_107_ ;
wire \IDU/Control/_108_ ;
wire \IDU/Control/_109_ ;
wire \IDU/Control/_110_ ;
wire \IDU/Control/_111_ ;
wire \IDU/Control/_112_ ;
wire \IDU/Control/_113_ ;
wire \IDU/Control/_114_ ;
wire \IDU/Control/_115_ ;
wire \IDU/Control/_116_ ;
wire \IDU/Control/_117_ ;
wire \IDU/Control/_118_ ;
wire \IDU/Control/_119_ ;
wire \IDU/Control/_120_ ;
wire \IDU/ImmGen/_000_ ;
wire \IDU/ImmGen/_001_ ;
wire \IDU/ImmGen/_002_ ;
wire \IDU/ImmGen/_003_ ;
wire \IDU/ImmGen/_004_ ;
wire \IDU/ImmGen/_005_ ;
wire \IDU/ImmGen/_006_ ;
wire \IDU/ImmGen/_007_ ;
wire \IDU/ImmGen/_008_ ;
wire \IDU/ImmGen/_009_ ;
wire \IDU/ImmGen/_010_ ;
wire \IDU/ImmGen/_011_ ;
wire \IDU/ImmGen/_012_ ;
wire \IDU/ImmGen/_013_ ;
wire \IDU/ImmGen/_014_ ;
wire \IDU/ImmGen/_015_ ;
wire \IDU/ImmGen/_016_ ;
wire \IDU/ImmGen/_017_ ;
wire \IDU/ImmGen/_018_ ;
wire \IDU/ImmGen/_019_ ;
wire \IDU/ImmGen/_020_ ;
wire \IDU/ImmGen/_021_ ;
wire \IDU/ImmGen/_022_ ;
wire \IDU/ImmGen/_023_ ;
wire \IDU/ImmGen/_024_ ;
wire \IDU/ImmGen/_025_ ;
wire \IDU/ImmGen/_026_ ;
wire \IDU/ImmGen/_027_ ;
wire \IDU/ImmGen/_028_ ;
wire \IDU/ImmGen/_029_ ;
wire \IDU/ImmGen/_030_ ;
wire \IDU/ImmGen/_031_ ;
wire \IDU/ImmGen/_032_ ;
wire \IDU/ImmGen/_033_ ;
wire \IDU/ImmGen/_034_ ;
wire \IDU/ImmGen/_035_ ;
wire \IDU/ImmGen/_036_ ;
wire \IDU/ImmGen/_037_ ;
wire \IDU/ImmGen/_038_ ;
wire \IDU/ImmGen/_039_ ;
wire \IDU/ImmGen/_040_ ;
wire \IDU/ImmGen/_041_ ;
wire \IDU/ImmGen/_042_ ;
wire \IDU/ImmGen/_043_ ;
wire \IDU/ImmGen/_044_ ;
wire \IDU/ImmGen/_045_ ;
wire \IDU/ImmGen/_046_ ;
wire \IDU/ImmGen/_047_ ;
wire \IDU/ImmGen/_048_ ;
wire \IDU/ImmGen/_049_ ;
wire \IDU/ImmGen/_050_ ;
wire \IDU/ImmGen/_051_ ;
wire \IDU/ImmGen/_052_ ;
wire \IDU/ImmGen/_053_ ;
wire \IDU/ImmGen/_054_ ;
wire \IDU/ImmGen/_055_ ;
wire \IDU/ImmGen/_056_ ;
wire \IDU/ImmGen/_057_ ;
wire \IDU/ImmGen/_058_ ;
wire \IDU/ImmGen/_059_ ;
wire \IDU/ImmGen/_060_ ;
wire \IDU/ImmGen/_061_ ;
wire \IDU/ImmGen/_062_ ;
wire \IDU/ImmGen/_063_ ;
wire \IDU/ImmGen/_064_ ;
wire \IDU/ImmGen/_065_ ;
wire \IDU/ImmGen/_066_ ;
wire \IDU/ImmGen/_067_ ;
wire \IDU/ImmGen/_068_ ;
wire \IDU/ImmGen/_069_ ;
wire \IDU/ImmGen/_070_ ;
wire \IDU/ImmGen/_071_ ;
wire \IDU/ImmGen/_072_ ;
wire \IDU/ImmGen/_073_ ;
wire \IDU/ImmGen/_074_ ;
wire \IDU/ImmGen/_075_ ;
wire \IDU/ImmGen/_076_ ;
wire \IDU/ImmGen/_077_ ;
wire \IDU/ImmGen/_078_ ;
wire \IDU/ImmGen/_079_ ;
wire \IDU/ImmGen/_080_ ;
wire \IDU/ImmGen/_081_ ;
wire \IDU/ImmGen/_082_ ;
wire \IDU/ImmGen/_083_ ;
wire \IDU/ImmGen/_084_ ;
wire \IDU/ImmGen/_085_ ;
wire \IDU/ImmGen/_086_ ;
wire \IDU/ImmGen/_087_ ;
wire \IDU/ImmGen/_088_ ;
wire \IDU/ImmGen/_089_ ;
wire \IFU/_000_ ;
wire \IFU/_001_ ;
wire \IFU/_002_ ;
wire \IFU/_003_ ;
wire \IFU/_004_ ;
wire \IFU/_005_ ;
wire \IFU/_006_ ;
wire \IFU/_007_ ;
wire \IFU/_008_ ;
wire \IFU/_009_ ;
wire \IFU/_010_ ;
wire \IFU/_011_ ;
wire \IFU/_012_ ;
wire \IFU/_013_ ;
wire \IFU/_014_ ;
wire \IFU/_015_ ;
wire \IFU/_016_ ;
wire \IFU/_017_ ;
wire \IFU/_018_ ;
wire \IFU/_019_ ;
wire \IFU/_020_ ;
wire \IFU/_021_ ;
wire \IFU/_022_ ;
wire \IFU/_023_ ;
wire \IFU/_024_ ;
wire \IFU/_025_ ;
wire \IFU/_026_ ;
wire \IFU/_027_ ;
wire \IFU/_028_ ;
wire \IFU/_029_ ;
wire \IFU/_030_ ;
wire \IFU/_031_ ;
wire \IFU/_032_ ;
wire \IFU/_033_ ;
wire \IFU/_034_ ;
wire \IFU/_035_ ;
wire \IFU/_036_ ;
wire \IFU/_037_ ;
wire \IFU/_038_ ;
wire \IFU/_039_ ;
wire \IFU/_040_ ;
wire \IFU/_041_ ;
wire \IFU/_042_ ;
wire \IFU/_043_ ;
wire \IFU/_044_ ;
wire \IFU/_045_ ;
wire \IFU/_046_ ;
wire \IFU/_047_ ;
wire \IFU/_048_ ;
wire \IFU/_049_ ;
wire \IFU/_050_ ;
wire \IFU/_051_ ;
wire \IFU/_052_ ;
wire \IFU/_053_ ;
wire \IFU/_054_ ;
wire \IFU/_055_ ;
wire \IFU/_056_ ;
wire \IFU/_057_ ;
wire \IFU/_058_ ;
wire \IFU/_059_ ;
wire \IFU/_060_ ;
wire \IFU/_061_ ;
wire \IFU/_062_ ;
wire \IFU/_063_ ;
wire \IFU/_064_ ;
wire \IFU/_065_ ;
wire \IFU/_066_ ;
wire \IFU/_067_ ;
wire \IFU/_068_ ;
wire \IFU/_069_ ;
wire \IFU/_070_ ;
wire \IFU/_071_ ;
wire \IFU/_072_ ;
wire \IFU/_073_ ;
wire \IFU/_074_ ;
wire \IFU/_075_ ;
wire \IFU/_076_ ;
wire \IFU/_077_ ;
wire \IFU/_078_ ;
wire \IFU/_079_ ;
wire \IFU/_080_ ;
wire \IFU/_081_ ;
wire \IFU/_082_ ;
wire \IFU/_083_ ;
wire \IFU/_084_ ;
wire \IFU/_085_ ;
wire \IFU/_086_ ;
wire \IFU/_087_ ;
wire \IFU/_088_ ;
wire \IFU/_089_ ;
wire \IFU/_090_ ;
wire \IFU/_091_ ;
wire \IFU/_092_ ;
wire \IFU/_093_ ;
wire \IFU/_094_ ;
wire \IFU/_095_ ;
wire \IFU/_096_ ;
wire \IFU/_097_ ;
wire \IFU/_098_ ;
wire \IFU/_099_ ;
wire \IFU/_100_ ;
wire \IFU/_101_ ;
wire \IFU/_102_ ;
wire \IFU/_103_ ;
wire \IFU/_104_ ;
wire \IFU/_105_ ;
wire \IFU/_106_ ;
wire \IFU/_107_ ;
wire \IFU/_108_ ;
wire \IFU/_109_ ;
wire \IFU/_110_ ;
wire \IFU/_111_ ;
wire \IFU/_112_ ;
wire \IFU/_113_ ;
wire \IFU/_114_ ;
wire \IFU/_115_ ;
wire \IFU/_116_ ;
wire \IFU/_117_ ;
wire \IFU/_118_ ;
wire \IFU/_119_ ;
wire \IFU/_120_ ;
wire \IFU/_121_ ;
wire \IFU/_122_ ;
wire \IFU/_123_ ;
wire \IFU/_124_ ;
wire \IFU/_125_ ;
wire \IFU/_126_ ;
wire \IFU/_127_ ;
wire \IFU/_128_ ;
wire \IFU/_129_ ;
wire \IFU/_130_ ;
wire \IFU/_131_ ;
wire \IFU/_132_ ;
wire \IFU/_133_ ;
wire \IFU/_134_ ;
wire \IFU/_135_ ;
wire \IFU/_136_ ;
wire \IFU/_137_ ;
wire \IFU/_138_ ;
wire \IFU/_139_ ;
wire \IFU/_140_ ;
wire \IFU/_141_ ;
wire \IFU/_142_ ;
wire \IFU/_143_ ;
wire \IFU/_144_ ;
wire \IFU/_145_ ;
wire \IFU/_146_ ;
wire \IFU/_147_ ;
wire \IFU/_148_ ;
wire \IFU/_149_ ;
wire \IFU/_150_ ;
wire \IFU/_151_ ;
wire \IFU/_152_ ;
wire \IFU/_153_ ;
wire \IFU/_154_ ;
wire \IFU/_155_ ;
wire \IFU/_156_ ;
wire \IFU/_157_ ;
wire \IFU/_158_ ;
wire \IFU/_159_ ;
wire \IFU/_160_ ;
wire \IFU/_161_ ;
wire \IFU/_162_ ;
wire \IFU/_163_ ;
wire \IFU/_164_ ;
wire \IFU/_165_ ;
wire \IFU/_166_ ;
wire \IFU/_167_ ;
wire \IFU/_168_ ;
wire \IFU/_169_ ;
wire \IFU/_170_ ;
wire \IFU/_171_ ;
wire \IFU/_172_ ;
wire \IFU/_173_ ;
wire \IFU/_174_ ;
wire \IFU/_175_ ;
wire \IFU/_176_ ;
wire \IFU/_177_ ;
wire \IFU/_178_ ;
wire \IFU/_179_ ;
wire \IFU/_180_ ;
wire \IFU/_181_ ;
wire \IFU/_182_ ;
wire \IFU/_183_ ;
wire \IFU/_184_ ;
wire \IFU/_185_ ;
wire \IFU/_186_ ;
wire \IFU/_187_ ;
wire \IFU/_188_ ;
wire \IFU/_189_ ;
wire \IFU/_190_ ;
wire \IFU/_191_ ;
wire \IFU/_192_ ;
wire \IFU/_193_ ;
wire \IFU/_194_ ;
wire \IFU/_195_ ;
wire \IFU/_196_ ;
wire \IFU/_197_ ;
wire \IFU/_198_ ;
wire \IFU/_199_ ;
wire \IFU/_200_ ;
wire \IFU/_201_ ;
wire \IFU/_202_ ;
wire \IFU/_203_ ;
wire \IFU/_204_ ;
wire \IFU/_205_ ;
wire \IFU/_206_ ;
wire \IFU/_207_ ;
wire \IFU/_208_ ;
wire \IFU/_209_ ;
wire \IFU/_210_ ;
wire \IFU/_211_ ;
wire \IFU/_212_ ;
wire \IFU/_213_ ;
wire \IFU/_214_ ;
wire \IFU/_215_ ;
wire \IFU/_216_ ;
wire \IFU/_217_ ;
wire \IFU/_218_ ;
wire \IFU/_219_ ;
wire \IFU/_220_ ;
wire \IFU/_221_ ;
wire \IFU/_222_ ;
wire \IFU/_223_ ;
wire \IFU/_224_ ;
wire \IFU/_225_ ;
wire \IFU/_226_ ;
wire \IFU/_227_ ;
wire \IFU/_228_ ;
wire \IFU/_229_ ;
wire \IFU/_230_ ;
wire \IFU/_231_ ;
wire \IFU/_232_ ;
wire \IFU/_233_ ;
wire \IFU/_234_ ;
wire \IFU/_235_ ;
wire \IFU/_236_ ;
wire \IFU/_237_ ;
wire \IFU/_238_ ;
wire \IFU/_239_ ;
wire \IFU/_240_ ;
wire \IFU/_241_ ;
wire \IFU/_242_ ;
wire \IFU/_243_ ;
wire \IFU/_244_ ;
wire \IFU/_245_ ;
wire \IFU/_246_ ;
wire \IFU/_247_ ;
wire \IFU/_248_ ;
wire \IFU/_249_ ;
wire \IFU/_250_ ;
wire \IFU/_251_ ;
wire \IFU/_252_ ;
wire \IFU/_253_ ;
wire \IFU/_254_ ;
wire \IFU/_255_ ;
wire \IFU/_256_ ;
wire \IFU/_257_ ;
wire \IFU/_258_ ;
wire \IFU/_259_ ;
wire \IFU/_260_ ;
wire \IFU/_261_ ;
wire \IFU/_262_ ;
wire \IFU/_263_ ;
wire \IFU/_264_ ;
wire \IFU/_265_ ;
wire \IFU/_266_ ;
wire \IFU/_267_ ;
wire \IFU/_268_ ;
wire \IFU/_269_ ;
wire \IFU/_270_ ;
wire \IFU/_271_ ;
wire \IFU/_272_ ;
wire \IFU/_273_ ;
wire \IFU/_274_ ;
wire \IFU/_275_ ;
wire \IFU/_276_ ;
wire \IFU/_277_ ;
wire \IFU/_278_ ;
wire \IFU/_279_ ;
wire \IFU/_280_ ;
wire \IFU/_281_ ;
wire \IFU/_282_ ;
wire \IFU/_283_ ;
wire \IFU/_284_ ;
wire \IFU/_285_ ;
wire \IFU/_286_ ;
wire \IFU/_287_ ;
wire \IFU/_288_ ;
wire \IFU/_289_ ;
wire \IFU/_290_ ;
wire \IFU/_291_ ;
wire \IFU/_292_ ;
wire \IFU/_293_ ;
wire \IFU/_294_ ;
wire \IFU/_295_ ;
wire \IFU/_296_ ;
wire \IFU/_297_ ;
wire \IFU/_298_ ;
wire \IFU/_299_ ;
wire \IFU/_300_ ;
wire \IFU/_301_ ;
wire \IFU/_302_ ;
wire \IFU/_303_ ;
wire \IFU/_304_ ;
wire \IFU/_305_ ;
wire \IFU/_306_ ;
wire \IFU/_307_ ;
wire \IFU/_308_ ;
wire \IFU/_309_ ;
wire \IFU/_310_ ;
wire \IFU/_311_ ;
wire \IFU/_312_ ;
wire \IFU/_313_ ;
wire \IFU/_314_ ;
wire \IFU/_315_ ;
wire \IFU/_316_ ;
wire \IFU/_317_ ;
wire \IFU/_318_ ;
wire \IFU/_319_ ;
wire \IFU/_320_ ;
wire \IFU/_321_ ;
wire \IFU/_322_ ;
wire \IFU/_323_ ;
wire \IFU/_324_ ;
wire \IFU/_325_ ;
wire \IFU/_326_ ;
wire \IFU/_327_ ;
wire \IFU/_328_ ;
wire \IFU/_329_ ;
wire \IFU/_330_ ;
wire \IFU/_331_ ;
wire \IFU/_332_ ;
wire \IFU/_333_ ;
wire \IFU/_334_ ;
wire \IFU/_335_ ;
wire \IFU/_336_ ;
wire \IFU/_337_ ;
wire \IFU/_338_ ;
wire \IFU/_339_ ;
wire \IFU/_340_ ;
wire \IFU/_341_ ;
wire \IFU/_342_ ;
wire \IFU/_343_ ;
wire \IFU/_344_ ;
wire \IFU/_345_ ;
wire \IFU/_346_ ;
wire \IFU/_347_ ;
wire \IFU/_348_ ;
wire \IFU/_349_ ;
wire \IFU/_350_ ;
wire \IFU/_351_ ;
wire \IFU/_352_ ;
wire \IFU/_353_ ;
wire \IFU/_354_ ;
wire \IFU/_355_ ;
wire \IFU/_356_ ;
wire \IFU/_357_ ;
wire \IFU/_358_ ;
wire \IFU/_359_ ;
wire \IFU/_360_ ;
wire \IFU/_361_ ;
wire \IFU/_362_ ;
wire \IFU/_363_ ;
wire \IFU/_364_ ;
wire \IFU/_365_ ;
wire \IFU/_366_ ;
wire \IFU/_367_ ;
wire \IFU/_368_ ;
wire \IFU/_369_ ;
wire \IFU/_370_ ;
wire \IFU/_371_ ;
wire \IFU/_372_ ;
wire \IFU/_373_ ;
wire \IFU/_374_ ;
wire \IFU/_375_ ;
wire \IFU/_376_ ;
wire \IFU/_377_ ;
wire \IFU/_378_ ;
wire \IFU/_379_ ;
wire \IFU/_380_ ;
wire \IFU/_381_ ;
wire \IFU/_382_ ;
wire \IFU/_383_ ;
wire \IFU/_384_ ;
wire \IFU/_385_ ;
wire \IFU/_386_ ;
wire \IFU/_387_ ;
wire \IFU/_388_ ;
wire \IFU/_389_ ;
wire \IFU/_390_ ;
wire \IFU/_391_ ;
wire \IFU/_392_ ;
wire \IFU/_393_ ;
wire \IFU/_394_ ;
wire \IFU/_395_ ;
wire \IFU/_396_ ;
wire \IFU/_397_ ;
wire \IFU/_398_ ;
wire \IFU/_399_ ;
wire \IFU/_400_ ;
wire \IFU/_401_ ;
wire \IFU/_402_ ;
wire \IFU/_403_ ;
wire \IFU/_404_ ;
wire \IFU/_405_ ;
wire \IFU/_406_ ;
wire \IFU/_407_ ;
wire \IFU/_408_ ;
wire \IFU/_409_ ;
wire \IFU/_410_ ;
wire \IFU/_411_ ;
wire \IFU/_412_ ;
wire \IFU/_413_ ;
wire \IFU/_414_ ;
wire \IFU/_415_ ;
wire \IFU/_416_ ;
wire \IFU/_417_ ;
wire \IFU/_418_ ;
wire \IFU/_419_ ;
wire \IFU/_420_ ;
wire \IFU/_421_ ;
wire \IFU/_422_ ;
wire \IFU/_423_ ;
wire \LSU/_0000_ ;
wire \LSU/_0001_ ;
wire \LSU/_0002_ ;
wire \LSU/_0003_ ;
wire \LSU/_0004_ ;
wire \LSU/_0005_ ;
wire \LSU/_0006_ ;
wire \LSU/_0007_ ;
wire \LSU/_0008_ ;
wire \LSU/_0009_ ;
wire \LSU/_0010_ ;
wire \LSU/_0011_ ;
wire \LSU/_0012_ ;
wire \LSU/_0013_ ;
wire \LSU/_0014_ ;
wire \LSU/_0015_ ;
wire \LSU/_0016_ ;
wire \LSU/_0017_ ;
wire \LSU/_0018_ ;
wire \LSU/_0019_ ;
wire \LSU/_0020_ ;
wire \LSU/_0021_ ;
wire \LSU/_0022_ ;
wire \LSU/_0023_ ;
wire \LSU/_0024_ ;
wire \LSU/_0025_ ;
wire \LSU/_0026_ ;
wire \LSU/_0027_ ;
wire \LSU/_0028_ ;
wire \LSU/_0029_ ;
wire \LSU/_0030_ ;
wire \LSU/_0031_ ;
wire \LSU/_0032_ ;
wire \LSU/_0033_ ;
wire \LSU/_0034_ ;
wire \LSU/_0035_ ;
wire \LSU/_0036_ ;
wire \LSU/_0037_ ;
wire \LSU/_0038_ ;
wire \LSU/_0039_ ;
wire \LSU/_0040_ ;
wire \LSU/_0041_ ;
wire \LSU/_0042_ ;
wire \LSU/_0043_ ;
wire \LSU/_0044_ ;
wire \LSU/_0045_ ;
wire \LSU/_0046_ ;
wire \LSU/_0047_ ;
wire \LSU/_0048_ ;
wire \LSU/_0049_ ;
wire \LSU/_0050_ ;
wire \LSU/_0051_ ;
wire \LSU/_0052_ ;
wire \LSU/_0053_ ;
wire \LSU/_0054_ ;
wire \LSU/_0055_ ;
wire \LSU/_0056_ ;
wire \LSU/_0057_ ;
wire \LSU/_0058_ ;
wire \LSU/_0059_ ;
wire \LSU/_0060_ ;
wire \LSU/_0061_ ;
wire \LSU/_0062_ ;
wire \LSU/_0063_ ;
wire \LSU/_0064_ ;
wire \LSU/_0065_ ;
wire \LSU/_0066_ ;
wire \LSU/_0067_ ;
wire \LSU/_0068_ ;
wire \LSU/_0069_ ;
wire \LSU/_0070_ ;
wire \LSU/_0071_ ;
wire \LSU/_0072_ ;
wire \LSU/_0073_ ;
wire \LSU/_0074_ ;
wire \LSU/_0075_ ;
wire \LSU/_0076_ ;
wire \LSU/_0077_ ;
wire \LSU/_0078_ ;
wire \LSU/_0079_ ;
wire \LSU/_0080_ ;
wire \LSU/_0081_ ;
wire \LSU/_0082_ ;
wire \LSU/_0083_ ;
wire \LSU/_0084_ ;
wire \LSU/_0085_ ;
wire \LSU/_0086_ ;
wire \LSU/_0087_ ;
wire \LSU/_0088_ ;
wire \LSU/_0089_ ;
wire \LSU/_0090_ ;
wire \LSU/_0091_ ;
wire \LSU/_0092_ ;
wire \LSU/_0093_ ;
wire \LSU/_0094_ ;
wire \LSU/_0095_ ;
wire \LSU/_0096_ ;
wire \LSU/_0097_ ;
wire \LSU/_0098_ ;
wire \LSU/_0099_ ;
wire \LSU/_0100_ ;
wire \LSU/_0101_ ;
wire \LSU/_0102_ ;
wire \LSU/_0103_ ;
wire \LSU/_0104_ ;
wire \LSU/_0105_ ;
wire \LSU/_0106_ ;
wire \LSU/_0107_ ;
wire \LSU/_0108_ ;
wire \LSU/_0109_ ;
wire \LSU/_0110_ ;
wire \LSU/_0111_ ;
wire \LSU/_0112_ ;
wire \LSU/_0113_ ;
wire \LSU/_0114_ ;
wire \LSU/_0115_ ;
wire \LSU/_0116_ ;
wire \LSU/_0117_ ;
wire \LSU/_0118_ ;
wire \LSU/_0119_ ;
wire \LSU/_0120_ ;
wire \LSU/_0121_ ;
wire \LSU/_0122_ ;
wire \LSU/_0123_ ;
wire \LSU/_0124_ ;
wire \LSU/_0125_ ;
wire \LSU/_0126_ ;
wire \LSU/_0127_ ;
wire \LSU/_0128_ ;
wire \LSU/_0129_ ;
wire \LSU/_0130_ ;
wire \LSU/_0131_ ;
wire \LSU/_0132_ ;
wire \LSU/_0133_ ;
wire \LSU/_0134_ ;
wire \LSU/_0135_ ;
wire \LSU/_0136_ ;
wire \LSU/_0137_ ;
wire \LSU/_0138_ ;
wire \LSU/_0139_ ;
wire \LSU/_0140_ ;
wire \LSU/_0141_ ;
wire \LSU/_0142_ ;
wire \LSU/_0143_ ;
wire \LSU/_0144_ ;
wire \LSU/_0145_ ;
wire \LSU/_0146_ ;
wire \LSU/_0147_ ;
wire \LSU/_0148_ ;
wire \LSU/_0149_ ;
wire \LSU/_0150_ ;
wire \LSU/_0151_ ;
wire \LSU/_0152_ ;
wire \LSU/_0153_ ;
wire \LSU/_0154_ ;
wire \LSU/_0155_ ;
wire \LSU/_0156_ ;
wire \LSU/_0157_ ;
wire \LSU/_0158_ ;
wire \LSU/_0159_ ;
wire \LSU/_0160_ ;
wire \LSU/_0161_ ;
wire \LSU/_0162_ ;
wire \LSU/_0163_ ;
wire \LSU/_0164_ ;
wire \LSU/_0165_ ;
wire \LSU/_0166_ ;
wire \LSU/_0167_ ;
wire \LSU/_0168_ ;
wire \LSU/_0169_ ;
wire \LSU/_0170_ ;
wire \LSU/_0171_ ;
wire \LSU/_0172_ ;
wire \LSU/_0173_ ;
wire \LSU/_0174_ ;
wire \LSU/_0175_ ;
wire \LSU/_0176_ ;
wire \LSU/_0177_ ;
wire \LSU/_0178_ ;
wire \LSU/_0179_ ;
wire \LSU/_0180_ ;
wire \LSU/_0181_ ;
wire \LSU/_0182_ ;
wire \LSU/_0183_ ;
wire \LSU/_0184_ ;
wire \LSU/_0185_ ;
wire \LSU/_0186_ ;
wire \LSU/_0187_ ;
wire \LSU/_0188_ ;
wire \LSU/_0189_ ;
wire \LSU/_0190_ ;
wire \LSU/_0191_ ;
wire \LSU/_0192_ ;
wire \LSU/_0193_ ;
wire \LSU/_0194_ ;
wire \LSU/_0195_ ;
wire \LSU/_0196_ ;
wire \LSU/_0197_ ;
wire \LSU/_0198_ ;
wire \LSU/_0199_ ;
wire \LSU/_0200_ ;
wire \LSU/_0201_ ;
wire \LSU/_0202_ ;
wire \LSU/_0203_ ;
wire \LSU/_0204_ ;
wire \LSU/_0205_ ;
wire \LSU/_0206_ ;
wire \LSU/_0207_ ;
wire \LSU/_0208_ ;
wire \LSU/_0209_ ;
wire \LSU/_0210_ ;
wire \LSU/_0211_ ;
wire \LSU/_0212_ ;
wire \LSU/_0213_ ;
wire \LSU/_0214_ ;
wire \LSU/_0215_ ;
wire \LSU/_0216_ ;
wire \LSU/_0217_ ;
wire \LSU/_0218_ ;
wire \LSU/_0219_ ;
wire \LSU/_0220_ ;
wire \LSU/_0221_ ;
wire \LSU/_0222_ ;
wire \LSU/_0223_ ;
wire \LSU/_0224_ ;
wire \LSU/_0225_ ;
wire \LSU/_0226_ ;
wire \LSU/_0227_ ;
wire \LSU/_0228_ ;
wire \LSU/_0229_ ;
wire \LSU/_0230_ ;
wire \LSU/_0231_ ;
wire \LSU/_0232_ ;
wire \LSU/_0233_ ;
wire \LSU/_0234_ ;
wire \LSU/_0235_ ;
wire \LSU/_0236_ ;
wire \LSU/_0237_ ;
wire \LSU/_0238_ ;
wire \LSU/_0239_ ;
wire \LSU/_0240_ ;
wire \LSU/_0241_ ;
wire \LSU/_0242_ ;
wire \LSU/_0243_ ;
wire \LSU/_0244_ ;
wire \LSU/_0245_ ;
wire \LSU/_0246_ ;
wire \LSU/_0247_ ;
wire \LSU/_0248_ ;
wire \LSU/_0249_ ;
wire \LSU/_0250_ ;
wire \LSU/_0251_ ;
wire \LSU/_0252_ ;
wire \LSU/_0253_ ;
wire \LSU/_0254_ ;
wire \LSU/_0255_ ;
wire \LSU/_0256_ ;
wire \LSU/_0257_ ;
wire \LSU/_0258_ ;
wire \LSU/_0259_ ;
wire \LSU/_0260_ ;
wire \LSU/_0261_ ;
wire \LSU/_0262_ ;
wire \LSU/_0263_ ;
wire \LSU/_0264_ ;
wire \LSU/_0265_ ;
wire \LSU/_0266_ ;
wire \LSU/_0267_ ;
wire \LSU/_0268_ ;
wire \LSU/_0269_ ;
wire \LSU/_0270_ ;
wire \LSU/_0271_ ;
wire \LSU/_0272_ ;
wire \LSU/_0273_ ;
wire \LSU/_0274_ ;
wire \LSU/_0275_ ;
wire \LSU/_0276_ ;
wire \LSU/_0277_ ;
wire \LSU/_0278_ ;
wire \LSU/_0279_ ;
wire \LSU/_0280_ ;
wire \LSU/_0281_ ;
wire \LSU/_0282_ ;
wire \LSU/_0283_ ;
wire \LSU/_0284_ ;
wire \LSU/_0285_ ;
wire \LSU/_0286_ ;
wire \LSU/_0287_ ;
wire \LSU/_0288_ ;
wire \LSU/_0289_ ;
wire \LSU/_0290_ ;
wire \LSU/_0291_ ;
wire \LSU/_0292_ ;
wire \LSU/_0293_ ;
wire \LSU/_0294_ ;
wire \LSU/_0295_ ;
wire \LSU/_0296_ ;
wire \LSU/_0297_ ;
wire \LSU/_0298_ ;
wire \LSU/_0299_ ;
wire \LSU/_0300_ ;
wire \LSU/_0301_ ;
wire \LSU/_0302_ ;
wire \LSU/_0303_ ;
wire \LSU/_0304_ ;
wire \LSU/_0305_ ;
wire \LSU/_0306_ ;
wire \LSU/_0307_ ;
wire \LSU/_0308_ ;
wire \LSU/_0309_ ;
wire \LSU/_0310_ ;
wire \LSU/_0311_ ;
wire \LSU/_0312_ ;
wire \LSU/_0313_ ;
wire \LSU/_0314_ ;
wire \LSU/_0315_ ;
wire \LSU/_0316_ ;
wire \LSU/_0317_ ;
wire \LSU/_0318_ ;
wire \LSU/_0319_ ;
wire \LSU/_0320_ ;
wire \LSU/_0321_ ;
wire \LSU/_0322_ ;
wire \LSU/_0323_ ;
wire \LSU/_0324_ ;
wire \LSU/_0325_ ;
wire \LSU/_0326_ ;
wire \LSU/_0327_ ;
wire \LSU/_0328_ ;
wire \LSU/_0329_ ;
wire \LSU/_0330_ ;
wire \LSU/_0331_ ;
wire \LSU/_0332_ ;
wire \LSU/_0333_ ;
wire \LSU/_0334_ ;
wire \LSU/_0335_ ;
wire \LSU/_0336_ ;
wire \LSU/_0337_ ;
wire \LSU/_0338_ ;
wire \LSU/_0339_ ;
wire \LSU/_0340_ ;
wire \LSU/_0341_ ;
wire \LSU/_0342_ ;
wire \LSU/_0343_ ;
wire \LSU/_0344_ ;
wire \LSU/_0345_ ;
wire \LSU/_0346_ ;
wire \LSU/_0347_ ;
wire \LSU/_0348_ ;
wire \LSU/_0349_ ;
wire \LSU/_0350_ ;
wire \LSU/_0351_ ;
wire \LSU/_0352_ ;
wire \LSU/_0353_ ;
wire \LSU/_0354_ ;
wire \LSU/_0355_ ;
wire \LSU/_0356_ ;
wire \LSU/_0357_ ;
wire \LSU/_0358_ ;
wire \LSU/_0359_ ;
wire \LSU/_0360_ ;
wire \LSU/_0361_ ;
wire \LSU/_0362_ ;
wire \LSU/_0363_ ;
wire \LSU/_0364_ ;
wire \LSU/_0365_ ;
wire \LSU/_0366_ ;
wire \LSU/_0367_ ;
wire \LSU/_0368_ ;
wire \LSU/_0369_ ;
wire \LSU/_0370_ ;
wire \LSU/_0371_ ;
wire \LSU/_0372_ ;
wire \LSU/_0373_ ;
wire \LSU/_0374_ ;
wire \LSU/_0375_ ;
wire \LSU/_0376_ ;
wire \LSU/_0377_ ;
wire \LSU/_0378_ ;
wire \LSU/_0379_ ;
wire \LSU/_0380_ ;
wire \LSU/_0381_ ;
wire \LSU/_0382_ ;
wire \LSU/_0383_ ;
wire \LSU/_0384_ ;
wire \LSU/_0385_ ;
wire \LSU/_0386_ ;
wire \LSU/_0387_ ;
wire \LSU/_0388_ ;
wire \LSU/_0389_ ;
wire \LSU/_0390_ ;
wire \LSU/_0391_ ;
wire \LSU/_0392_ ;
wire \LSU/_0393_ ;
wire \LSU/_0394_ ;
wire \LSU/_0395_ ;
wire \LSU/_0396_ ;
wire \LSU/_0397_ ;
wire \LSU/_0398_ ;
wire \LSU/_0399_ ;
wire \LSU/_0400_ ;
wire \LSU/_0401_ ;
wire \LSU/_0402_ ;
wire \LSU/_0403_ ;
wire \LSU/_0404_ ;
wire \LSU/_0405_ ;
wire \LSU/_0406_ ;
wire \LSU/_0407_ ;
wire \LSU/_0408_ ;
wire \LSU/_0409_ ;
wire \LSU/_0410_ ;
wire \LSU/_0411_ ;
wire \LSU/_0412_ ;
wire \LSU/_0413_ ;
wire \LSU/_0414_ ;
wire \LSU/_0415_ ;
wire \LSU/_0416_ ;
wire \LSU/_0417_ ;
wire \LSU/_0418_ ;
wire \LSU/_0419_ ;
wire \LSU/_0420_ ;
wire \LSU/_0421_ ;
wire \LSU/_0422_ ;
wire \LSU/_0423_ ;
wire \LSU/_0424_ ;
wire \LSU/_0425_ ;
wire \LSU/_0426_ ;
wire \LSU/_0427_ ;
wire \LSU/_0428_ ;
wire \LSU/_0429_ ;
wire \LSU/_0430_ ;
wire \LSU/_0431_ ;
wire \LSU/_0432_ ;
wire \LSU/_0433_ ;
wire \LSU/_0434_ ;
wire \LSU/_0435_ ;
wire \LSU/_0436_ ;
wire \LSU/_0437_ ;
wire \LSU/_0438_ ;
wire \LSU/_0439_ ;
wire \LSU/_0440_ ;
wire \LSU/_0441_ ;
wire \LSU/_0442_ ;
wire \LSU/_0443_ ;
wire \LSU/_0444_ ;
wire \LSU/_0445_ ;
wire \LSU/_0446_ ;
wire \LSU/_0447_ ;
wire \LSU/_0448_ ;
wire \LSU/_0449_ ;
wire \LSU/_0450_ ;
wire \LSU/_0451_ ;
wire \LSU/_0452_ ;
wire \LSU/_0453_ ;
wire \LSU/_0454_ ;
wire \LSU/_0455_ ;
wire \LSU/_0456_ ;
wire \LSU/_0457_ ;
wire \LSU/_0458_ ;
wire \LSU/_0459_ ;
wire \LSU/_0460_ ;
wire \LSU/_0461_ ;
wire \LSU/_0462_ ;
wire \LSU/_0463_ ;
wire \LSU/_0464_ ;
wire \LSU/_0465_ ;
wire \LSU/_0466_ ;
wire \LSU/_0467_ ;
wire \LSU/_0468_ ;
wire \LSU/_0469_ ;
wire \LSU/_0470_ ;
wire \LSU/_0471_ ;
wire \LSU/_0472_ ;
wire \LSU/_0473_ ;
wire \LSU/_0474_ ;
wire \LSU/_0475_ ;
wire \LSU/_0476_ ;
wire \LSU/_0477_ ;
wire \LSU/_0478_ ;
wire \LSU/_0479_ ;
wire \LSU/_0480_ ;
wire \LSU/_0481_ ;
wire \LSU/_0482_ ;
wire \LSU/_0483_ ;
wire \LSU/_0484_ ;
wire \LSU/_0485_ ;
wire \LSU/_0486_ ;
wire \LSU/_0487_ ;
wire \LSU/_0488_ ;
wire \LSU/_0489_ ;
wire \LSU/_0490_ ;
wire \LSU/_0491_ ;
wire \LSU/_0492_ ;
wire \LSU/_0493_ ;
wire \LSU/_0494_ ;
wire \LSU/_0495_ ;
wire \LSU/_0496_ ;
wire \LSU/_0497_ ;
wire \LSU/_0498_ ;
wire \LSU/_0499_ ;
wire \LSU/_0500_ ;
wire \LSU/_0501_ ;
wire \LSU/_0502_ ;
wire \LSU/_0503_ ;
wire \LSU/_0504_ ;
wire \LSU/_0505_ ;
wire \LSU/_0506_ ;
wire \LSU/_0507_ ;
wire \LSU/_0508_ ;
wire \LSU/_0509_ ;
wire \LSU/_0510_ ;
wire \LSU/_0511_ ;
wire \LSU/_0512_ ;
wire \LSU/_0513_ ;
wire \LSU/_0514_ ;
wire \LSU/_0515_ ;
wire \LSU/_0516_ ;
wire \LSU/_0517_ ;
wire \LSU/_0518_ ;
wire \LSU/_0519_ ;
wire \LSU/_0520_ ;
wire \LSU/_0521_ ;
wire \LSU/_0522_ ;
wire \LSU/_0523_ ;
wire \LSU/_0524_ ;
wire \LSU/_0525_ ;
wire \LSU/_0526_ ;
wire \LSU/_0527_ ;
wire \LSU/_0528_ ;
wire \LSU/_0529_ ;
wire \LSU/_0530_ ;
wire \LSU/_0531_ ;
wire \LSU/_0532_ ;
wire \LSU/_0533_ ;
wire \LSU/_0534_ ;
wire \LSU/_0535_ ;
wire \LSU/_0536_ ;
wire \LSU/_0537_ ;
wire \LSU/_0538_ ;
wire \LSU/_0539_ ;
wire \LSU/_0540_ ;
wire \LSU/_0541_ ;
wire \LSU/_0542_ ;
wire \LSU/_0543_ ;
wire \LSU/_0544_ ;
wire \LSU/_0545_ ;
wire \LSU/_0546_ ;
wire \LSU/_0547_ ;
wire \LSU/_0548_ ;
wire \LSU/_0549_ ;
wire \LSU/_0550_ ;
wire \LSU/_0551_ ;
wire \LSU/_0552_ ;
wire \LSU/_0553_ ;
wire \LSU/_0554_ ;
wire \LSU/_0555_ ;
wire \LSU/_0556_ ;
wire \LSU/_0557_ ;
wire \LSU/_0558_ ;
wire \LSU/_0559_ ;
wire \LSU/_0560_ ;
wire \LSU/_0561_ ;
wire \LSU/_0562_ ;
wire \LSU/_0563_ ;
wire \LSU/_0564_ ;
wire \LSU/_0565_ ;
wire \LSU/_0566_ ;
wire \LSU/_0567_ ;
wire \LSU/_0568_ ;
wire \LSU/_0569_ ;
wire \LSU/_0570_ ;
wire \LSU/_0571_ ;
wire \LSU/_0572_ ;
wire \LSU/_0573_ ;
wire \LSU/_0574_ ;
wire \LSU/_0575_ ;
wire \LSU/_0576_ ;
wire \LSU/_0577_ ;
wire \LSU/_0578_ ;
wire \LSU/_0579_ ;
wire \LSU/_0580_ ;
wire \LSU/_0581_ ;
wire \LSU/_0582_ ;
wire \LSU/_0583_ ;
wire \LSU/_0584_ ;
wire \LSU/_0585_ ;
wire \LSU/_0586_ ;
wire \LSU/_0587_ ;
wire \LSU/_0588_ ;
wire \LSU/_0589_ ;
wire \LSU/_0590_ ;
wire \LSU/_0591_ ;
wire \LSU/_0592_ ;
wire \LSU/_0593_ ;
wire \LSU/_0594_ ;
wire \LSU/_0595_ ;
wire \LSU/_0596_ ;
wire \LSU/_0597_ ;
wire \LSU/_0598_ ;
wire \LSU/_0599_ ;
wire \LSU/_0600_ ;
wire \LSU/_0601_ ;
wire \LSU/_0602_ ;
wire \LSU/_0603_ ;
wire \LSU/_0604_ ;
wire \LSU/_0605_ ;
wire \LSU/_0606_ ;
wire \LSU/_0607_ ;
wire \LSU/_0608_ ;
wire \LSU/_0609_ ;
wire \LSU/_0610_ ;
wire \LSU/_0611_ ;
wire \LSU/_0612_ ;
wire \LSU/_0613_ ;
wire \LSU/_0614_ ;
wire \LSU/_0615_ ;
wire \LSU/_0616_ ;
wire \LSU/_0617_ ;
wire \LSU/_0618_ ;
wire \LSU/_0619_ ;
wire \LSU/_0620_ ;
wire \LSU/_0621_ ;
wire \LSU/_0622_ ;
wire \LSU/_0623_ ;
wire \LSU/_0624_ ;
wire \LSU/_0625_ ;
wire \LSU/_0626_ ;
wire \LSU/_0627_ ;
wire \LSU/_0628_ ;
wire \LSU/_0629_ ;
wire \LSU/_0630_ ;
wire \LSU/_0631_ ;
wire \LSU/_0632_ ;
wire \LSU/_0633_ ;
wire \LSU/_0634_ ;
wire \LSU/_0635_ ;
wire \LSU/_0636_ ;
wire \LSU/_0637_ ;
wire \LSU/_0638_ ;
wire \LSU/_0639_ ;
wire \LSU/_0640_ ;
wire \LSU/_0641_ ;
wire \LSU/_0642_ ;
wire \LSU/_0643_ ;
wire \LSU/_0644_ ;
wire \LSU/_0645_ ;
wire \LSU/_0646_ ;
wire \LSU/_0647_ ;
wire \LSU/_0648_ ;
wire \LSU/_0649_ ;
wire \LSU/_0650_ ;
wire \LSU/_0651_ ;
wire \LSU/_0652_ ;
wire \LSU/_0653_ ;
wire \LSU/_0654_ ;
wire \LSU/_0655_ ;
wire \LSU/_0656_ ;
wire \LSU/_0657_ ;
wire \LSU/_0658_ ;
wire \LSU/_0659_ ;
wire \LSU/_0660_ ;
wire \LSU/_0661_ ;
wire \LSU/_0662_ ;
wire \LSU/_0663_ ;
wire \LSU/_0664_ ;
wire \LSU/_0665_ ;
wire \LSU/_0666_ ;
wire \LSU/_0667_ ;
wire \LSU/_0668_ ;
wire \LSU/_0669_ ;
wire \LSU/_0670_ ;
wire \LSU/_0671_ ;
wire \LSU/_0672_ ;
wire \LSU/_0673_ ;
wire \LSU/_0674_ ;
wire \LSU/_0675_ ;
wire \LSU/_0676_ ;
wire \LSU/_0677_ ;
wire \LSU/_0678_ ;
wire \LSU/_0679_ ;
wire \LSU/_0680_ ;
wire \LSU/_0681_ ;
wire \LSU/_0682_ ;
wire \LSU/_0683_ ;
wire \LSU/_0684_ ;
wire \LSU/_0685_ ;
wire \LSU/_0686_ ;
wire \LSU/_0687_ ;
wire \LSU/_0688_ ;
wire \LSU/_0689_ ;
wire \LSU/_0690_ ;
wire \LSU/_0691_ ;
wire \LSU/_0692_ ;
wire \LSU/_0693_ ;
wire \LSU/_0694_ ;
wire \LSU/_0695_ ;
wire \LSU/_0696_ ;
wire \LSU/_0697_ ;
wire \LSU/_0698_ ;
wire \LSU/_0699_ ;
wire \LSU/_0700_ ;
wire \LSU/_0701_ ;
wire \LSU/_0702_ ;
wire \LSU/_0703_ ;
wire \LSU/_0704_ ;
wire \LSU/_0705_ ;
wire \LSU/_0706_ ;
wire \LSU/_0707_ ;
wire \LSU/_0708_ ;
wire \LSU/_0709_ ;
wire \LSU/_0710_ ;
wire \LSU/_0711_ ;
wire \LSU/_0712_ ;
wire \LSU/_0713_ ;
wire \LSU/_0714_ ;
wire \LSU/_0715_ ;
wire \LSU/_0716_ ;
wire \LSU/_0717_ ;
wire \LSU/_0718_ ;
wire \LSU/_0719_ ;
wire \LSU/_0720_ ;
wire \LSU/_0721_ ;
wire \LSU/_0722_ ;
wire \LSU/_0723_ ;
wire \LSU/_0724_ ;
wire \LSU/_0725_ ;
wire \LSU/_0726_ ;
wire \LSU/_0727_ ;
wire \LSU/_0728_ ;
wire \LSU/_0729_ ;
wire \LSU/_0730_ ;
wire \LSU/_0731_ ;
wire \LSU/_0732_ ;
wire \LSU/_0733_ ;
wire \LSU/_0734_ ;
wire \LSU/_0735_ ;
wire \LSU/_0736_ ;
wire \LSU/_0737_ ;
wire \LSU/_0738_ ;
wire \LSU/_0739_ ;
wire \LSU/_0740_ ;
wire \LSU/_0741_ ;
wire \LSU/_0742_ ;
wire \LSU/_0743_ ;
wire \LSU/_0744_ ;
wire \LSU/_0745_ ;
wire \LSU/_0746_ ;
wire \LSU/_0747_ ;
wire \LSU/_0748_ ;
wire \LSU/_0749_ ;
wire \LSU/_0750_ ;
wire \LSU/_0751_ ;
wire \LSU/_0752_ ;
wire \LSU/_0753_ ;
wire \LSU/_0754_ ;
wire \LSU/_0755_ ;
wire \LSU/_0756_ ;
wire \LSU/_0757_ ;
wire \LSU/_0758_ ;
wire \LSU/_0759_ ;
wire \LSU/_0760_ ;
wire \LSU/_0761_ ;
wire \LSU/_0762_ ;
wire \LSU/_0763_ ;
wire \LSU/_0764_ ;
wire \LSU/_0765_ ;
wire \LSU/_0766_ ;
wire \LSU/_0767_ ;
wire \LSU/_0768_ ;
wire \LSU/_0769_ ;
wire \LSU/_0770_ ;
wire \LSU/_0771_ ;
wire \LSU/_0772_ ;
wire \LSU/_0773_ ;
wire \LSU/_0774_ ;
wire \LSU/_0775_ ;
wire \LSU/_0776_ ;
wire \LSU/_0777_ ;
wire \LSU/_0778_ ;
wire \LSU/_0779_ ;
wire \LSU/_0780_ ;
wire \LSU/_0781_ ;
wire \LSU/_0782_ ;
wire \LSU/_0783_ ;
wire \LSU/_0784_ ;
wire \LSU/_0785_ ;
wire \LSU/_0786_ ;
wire \LSU/_0787_ ;
wire \LSU/_0788_ ;
wire \LSU/_0789_ ;
wire \LSU/_0790_ ;
wire \LSU/_0791_ ;
wire \LSU/_0792_ ;
wire \LSU/_0793_ ;
wire \LSU/_0794_ ;
wire \LSU/_0795_ ;
wire \LSU/_0796_ ;
wire \LSU/_0797_ ;
wire \LSU/_0798_ ;
wire \LSU/_0799_ ;
wire \LSU/_0800_ ;
wire \LSU/_0801_ ;
wire \LSU/_0802_ ;
wire \LSU/_0803_ ;
wire \LSU/_0804_ ;
wire \LSU/_0805_ ;
wire \LSU/_0806_ ;
wire \LSU/_0807_ ;
wire \LSU/_0808_ ;
wire \LSU/_0809_ ;
wire \LSU/_0810_ ;
wire \LSU/_0811_ ;
wire \LSU/_0812_ ;
wire \LSU/_0813_ ;
wire \LSU/_0814_ ;
wire \LSU/_0815_ ;
wire \LSU/_0816_ ;
wire \LSU/_0817_ ;
wire \LSU/_0818_ ;
wire \LSU/_0819_ ;
wire \LSU/_0820_ ;
wire \LSU/_0821_ ;
wire \LSU/_0822_ ;
wire \LSU/_0823_ ;
wire \LSU/_0824_ ;
wire \LSU/_0825_ ;
wire \LSU/_0826_ ;
wire \LSU/_0827_ ;
wire \LSU/_0828_ ;
wire \LSU/_0829_ ;
wire \LSU/_0830_ ;
wire \LSU/_0831_ ;
wire \LSU/_0832_ ;
wire \LSU/_0833_ ;
wire \LSU/_0834_ ;
wire \LSU/_0835_ ;
wire \LSU/_0836_ ;
wire \LSU/_0837_ ;
wire \LSU/_0838_ ;
wire \LSU/_0839_ ;
wire \LSU/_0840_ ;
wire \LSU/_0841_ ;
wire \LSU/_0842_ ;
wire \LSU/_0843_ ;
wire \LSU/_0844_ ;
wire \LSU/_0845_ ;
wire \LSU/_0846_ ;
wire \LSU/_0847_ ;
wire \LSU/_0848_ ;
wire \LSU/_0849_ ;
wire \LSU/_0850_ ;
wire \LSU/_0851_ ;
wire \LSU/_0852_ ;
wire \LSU/_0853_ ;
wire \LSU/_0854_ ;
wire \LSU/_0855_ ;
wire \LSU/_0856_ ;
wire \LSU/_0857_ ;
wire \LSU/_0858_ ;
wire \LSU/_0859_ ;
wire \LSU/_0860_ ;
wire \LSU/_0861_ ;
wire \LSU/_0862_ ;
wire \LSU/_0863_ ;
wire \LSU/_0864_ ;
wire \LSU/_0865_ ;
wire \LSU/_0866_ ;
wire \LSU/_0867_ ;
wire \LSU/_0868_ ;
wire \LSU/_0869_ ;
wire \LSU/_0870_ ;
wire \LSU/_0871_ ;
wire \LSU/_0872_ ;
wire \LSU/_0873_ ;
wire \LSU/_0874_ ;
wire \LSU/_0875_ ;
wire \LSU/_0876_ ;
wire \LSU/_0877_ ;
wire \LSU/_0878_ ;
wire \LSU/_0879_ ;
wire \LSU/_0880_ ;
wire \LSU/_0881_ ;
wire \LSU/_0882_ ;
wire \LSU/_0883_ ;
wire \LSU/_0884_ ;
wire \LSU/_0885_ ;
wire \LSU/_0886_ ;
wire \LSU/_0887_ ;
wire \LSU/_0888_ ;
wire \LSU/_0889_ ;
wire \LSU/_0890_ ;
wire \LSU/_0891_ ;
wire \LSU/_0892_ ;
wire \LSU/_0893_ ;
wire \LSU/_0894_ ;
wire \LSU/_0895_ ;
wire \LSU/_0896_ ;
wire \LSU/_0897_ ;
wire \LSU/_0898_ ;
wire \LSU/_0899_ ;
wire \LSU/_0900_ ;
wire \LSU/_0901_ ;
wire \LSU/_0902_ ;
wire \LSU/_0903_ ;
wire \LSU/_0904_ ;
wire \LSU/_0905_ ;
wire \LSU/_0906_ ;
wire \LSU/_0907_ ;
wire \LSU/_0908_ ;
wire \LSU/_0909_ ;
wire \LSU/_0910_ ;
wire \LSU/_0911_ ;
wire \LSU/_0912_ ;
wire \LSU/_0913_ ;
wire \LSU/_0914_ ;
wire \LSU/_0915_ ;
wire \LSU/_0916_ ;
wire \LSU/_0917_ ;
wire \LSU/_0918_ ;
wire \LSU/_0919_ ;
wire \LSU/_0920_ ;
wire \LSU/_0921_ ;
wire \LSU/_0922_ ;
wire \LSU/_0923_ ;
wire \LSU/_0924_ ;
wire \LSU/_0925_ ;
wire \LSU/_0926_ ;
wire \LSU/_0927_ ;
wire \LSU/_0928_ ;
wire \LSU/_0929_ ;
wire \LSU/_0930_ ;
wire \LSU/_0931_ ;
wire \LSU/_0932_ ;
wire \LSU/_0933_ ;
wire \LSU/_0934_ ;
wire \LSU/_0935_ ;
wire \LSU/_0936_ ;
wire \LSU/_0937_ ;
wire \LSU/_0938_ ;
wire \LSU/_0939_ ;
wire \LSU/_0940_ ;
wire \LSU/_0941_ ;
wire \LSU/_0942_ ;
wire \LSU/_0943_ ;
wire \LSU/_0944_ ;
wire \LSU/_0945_ ;
wire \LSU/_0946_ ;
wire \LSU/_0947_ ;
wire \LSU/_0948_ ;
wire \LSU/_0949_ ;
wire \LSU/_0950_ ;
wire \LSU/_0951_ ;
wire \LSU/_0952_ ;
wire \LSU/_0953_ ;
wire \LSU/_0954_ ;
wire \LSU/_0955_ ;
wire \LSU/_0956_ ;
wire \LSU/_0957_ ;
wire \LSU/_0958_ ;
wire \LSU/_0959_ ;
wire \LSU/_0960_ ;
wire \LSU/_0961_ ;
wire \LSU/_0962_ ;
wire \LSU/_0963_ ;
wire \LSU/_0964_ ;
wire \LSU/_0965_ ;
wire \LSU/_0966_ ;
wire \LSU/_0967_ ;
wire \LSU/_0968_ ;
wire \LSU/_0969_ ;
wire \LSU/_0970_ ;
wire \LSU/_0971_ ;
wire \LSU/_0972_ ;
wire \LSU/_0973_ ;
wire \LSU/_0974_ ;
wire \LSU/_0975_ ;
wire \LSU/_0976_ ;
wire \LSU/_0977_ ;
wire \LSU/_0978_ ;
wire \LSU/_0979_ ;
wire \LSU/_0980_ ;
wire \LSU/_0981_ ;
wire \LSU/_0982_ ;
wire \LSU/_0983_ ;
wire \RegFile/_0000_ ;
wire \RegFile/_0001_ ;
wire \RegFile/_0002_ ;
wire \RegFile/_0003_ ;
wire \RegFile/_0004_ ;
wire \RegFile/_0005_ ;
wire \RegFile/_0006_ ;
wire \RegFile/_0007_ ;
wire \RegFile/_0008_ ;
wire \RegFile/_0009_ ;
wire \RegFile/_0010_ ;
wire \RegFile/_0011_ ;
wire \RegFile/_0012_ ;
wire \RegFile/_0013_ ;
wire \RegFile/_0014_ ;
wire \RegFile/_0015_ ;
wire \RegFile/_0016_ ;
wire \RegFile/_0017_ ;
wire \RegFile/_0018_ ;
wire \RegFile/_0019_ ;
wire \RegFile/_0020_ ;
wire \RegFile/_0021_ ;
wire \RegFile/_0022_ ;
wire \RegFile/_0023_ ;
wire \RegFile/_0024_ ;
wire \RegFile/_0025_ ;
wire \RegFile/_0026_ ;
wire \RegFile/_0027_ ;
wire \RegFile/_0028_ ;
wire \RegFile/_0029_ ;
wire \RegFile/_0030_ ;
wire \RegFile/_0031_ ;
wire \RegFile/_0032_ ;
wire \RegFile/_0033_ ;
wire \RegFile/_0034_ ;
wire \RegFile/_0035_ ;
wire \RegFile/_0036_ ;
wire \RegFile/_0037_ ;
wire \RegFile/_0038_ ;
wire \RegFile/_0039_ ;
wire \RegFile/_0040_ ;
wire \RegFile/_0041_ ;
wire \RegFile/_0042_ ;
wire \RegFile/_0043_ ;
wire \RegFile/_0044_ ;
wire \RegFile/_0045_ ;
wire \RegFile/_0046_ ;
wire \RegFile/_0047_ ;
wire \RegFile/_0048_ ;
wire \RegFile/_0049_ ;
wire \RegFile/_0050_ ;
wire \RegFile/_0051_ ;
wire \RegFile/_0052_ ;
wire \RegFile/_0053_ ;
wire \RegFile/_0054_ ;
wire \RegFile/_0055_ ;
wire \RegFile/_0056_ ;
wire \RegFile/_0057_ ;
wire \RegFile/_0058_ ;
wire \RegFile/_0059_ ;
wire \RegFile/_0060_ ;
wire \RegFile/_0061_ ;
wire \RegFile/_0062_ ;
wire \RegFile/_0063_ ;
wire \RegFile/_0064_ ;
wire \RegFile/_0065_ ;
wire \RegFile/_0066_ ;
wire \RegFile/_0067_ ;
wire \RegFile/_0068_ ;
wire \RegFile/_0069_ ;
wire \RegFile/_0070_ ;
wire \RegFile/_0071_ ;
wire \RegFile/_0072_ ;
wire \RegFile/_0073_ ;
wire \RegFile/_0074_ ;
wire \RegFile/_0075_ ;
wire \RegFile/_0076_ ;
wire \RegFile/_0077_ ;
wire \RegFile/_0078_ ;
wire \RegFile/_0079_ ;
wire \RegFile/_0080_ ;
wire \RegFile/_0081_ ;
wire \RegFile/_0082_ ;
wire \RegFile/_0083_ ;
wire \RegFile/_0084_ ;
wire \RegFile/_0085_ ;
wire \RegFile/_0086_ ;
wire \RegFile/_0087_ ;
wire \RegFile/_0088_ ;
wire \RegFile/_0089_ ;
wire \RegFile/_0090_ ;
wire \RegFile/_0091_ ;
wire \RegFile/_0092_ ;
wire \RegFile/_0093_ ;
wire \RegFile/_0094_ ;
wire \RegFile/_0095_ ;
wire \RegFile/_0096_ ;
wire \RegFile/_0097_ ;
wire \RegFile/_0098_ ;
wire \RegFile/_0099_ ;
wire \RegFile/_0100_ ;
wire \RegFile/_0101_ ;
wire \RegFile/_0102_ ;
wire \RegFile/_0103_ ;
wire \RegFile/_0104_ ;
wire \RegFile/_0105_ ;
wire \RegFile/_0106_ ;
wire \RegFile/_0107_ ;
wire \RegFile/_0108_ ;
wire \RegFile/_0109_ ;
wire \RegFile/_0110_ ;
wire \RegFile/_0111_ ;
wire \RegFile/_0112_ ;
wire \RegFile/_0113_ ;
wire \RegFile/_0114_ ;
wire \RegFile/_0115_ ;
wire \RegFile/_0116_ ;
wire \RegFile/_0117_ ;
wire \RegFile/_0118_ ;
wire \RegFile/_0119_ ;
wire \RegFile/_0120_ ;
wire \RegFile/_0121_ ;
wire \RegFile/_0122_ ;
wire \RegFile/_0123_ ;
wire \RegFile/_0124_ ;
wire \RegFile/_0125_ ;
wire \RegFile/_0126_ ;
wire \RegFile/_0127_ ;
wire \RegFile/_0128_ ;
wire \RegFile/_0129_ ;
wire \RegFile/_0130_ ;
wire \RegFile/_0131_ ;
wire \RegFile/_0132_ ;
wire \RegFile/_0133_ ;
wire \RegFile/_0134_ ;
wire \RegFile/_0135_ ;
wire \RegFile/_0136_ ;
wire \RegFile/_0137_ ;
wire \RegFile/_0138_ ;
wire \RegFile/_0139_ ;
wire \RegFile/_0140_ ;
wire \RegFile/_0141_ ;
wire \RegFile/_0142_ ;
wire \RegFile/_0143_ ;
wire \RegFile/_0144_ ;
wire \RegFile/_0145_ ;
wire \RegFile/_0146_ ;
wire \RegFile/_0147_ ;
wire \RegFile/_0148_ ;
wire \RegFile/_0149_ ;
wire \RegFile/_0150_ ;
wire \RegFile/_0151_ ;
wire \RegFile/_0152_ ;
wire \RegFile/_0153_ ;
wire \RegFile/_0154_ ;
wire \RegFile/_0155_ ;
wire \RegFile/_0156_ ;
wire \RegFile/_0157_ ;
wire \RegFile/_0158_ ;
wire \RegFile/_0159_ ;
wire \RegFile/_0160_ ;
wire \RegFile/_0161_ ;
wire \RegFile/_0162_ ;
wire \RegFile/_0163_ ;
wire \RegFile/_0164_ ;
wire \RegFile/_0165_ ;
wire \RegFile/_0166_ ;
wire \RegFile/_0167_ ;
wire \RegFile/_0168_ ;
wire \RegFile/_0169_ ;
wire \RegFile/_0170_ ;
wire \RegFile/_0171_ ;
wire \RegFile/_0172_ ;
wire \RegFile/_0173_ ;
wire \RegFile/_0174_ ;
wire \RegFile/_0175_ ;
wire \RegFile/_0176_ ;
wire \RegFile/_0177_ ;
wire \RegFile/_0178_ ;
wire \RegFile/_0179_ ;
wire \RegFile/_0180_ ;
wire \RegFile/_0181_ ;
wire \RegFile/_0182_ ;
wire \RegFile/_0183_ ;
wire \RegFile/_0184_ ;
wire \RegFile/_0185_ ;
wire \RegFile/_0186_ ;
wire \RegFile/_0187_ ;
wire \RegFile/_0188_ ;
wire \RegFile/_0189_ ;
wire \RegFile/_0190_ ;
wire \RegFile/_0191_ ;
wire \RegFile/_0192_ ;
wire \RegFile/_0193_ ;
wire \RegFile/_0194_ ;
wire \RegFile/_0195_ ;
wire \RegFile/_0196_ ;
wire \RegFile/_0197_ ;
wire \RegFile/_0198_ ;
wire \RegFile/_0199_ ;
wire \RegFile/_0200_ ;
wire \RegFile/_0201_ ;
wire \RegFile/_0202_ ;
wire \RegFile/_0203_ ;
wire \RegFile/_0204_ ;
wire \RegFile/_0205_ ;
wire \RegFile/_0206_ ;
wire \RegFile/_0207_ ;
wire \RegFile/_0208_ ;
wire \RegFile/_0209_ ;
wire \RegFile/_0210_ ;
wire \RegFile/_0211_ ;
wire \RegFile/_0212_ ;
wire \RegFile/_0213_ ;
wire \RegFile/_0214_ ;
wire \RegFile/_0215_ ;
wire \RegFile/_0216_ ;
wire \RegFile/_0217_ ;
wire \RegFile/_0218_ ;
wire \RegFile/_0219_ ;
wire \RegFile/_0220_ ;
wire \RegFile/_0221_ ;
wire \RegFile/_0222_ ;
wire \RegFile/_0223_ ;
wire \RegFile/_0224_ ;
wire \RegFile/_0225_ ;
wire \RegFile/_0226_ ;
wire \RegFile/_0227_ ;
wire \RegFile/_0228_ ;
wire \RegFile/_0229_ ;
wire \RegFile/_0230_ ;
wire \RegFile/_0231_ ;
wire \RegFile/_0232_ ;
wire \RegFile/_0233_ ;
wire \RegFile/_0234_ ;
wire \RegFile/_0235_ ;
wire \RegFile/_0236_ ;
wire \RegFile/_0237_ ;
wire \RegFile/_0238_ ;
wire \RegFile/_0239_ ;
wire \RegFile/_0240_ ;
wire \RegFile/_0241_ ;
wire \RegFile/_0242_ ;
wire \RegFile/_0243_ ;
wire \RegFile/_0244_ ;
wire \RegFile/_0245_ ;
wire \RegFile/_0246_ ;
wire \RegFile/_0247_ ;
wire \RegFile/_0248_ ;
wire \RegFile/_0249_ ;
wire \RegFile/_0250_ ;
wire \RegFile/_0251_ ;
wire \RegFile/_0252_ ;
wire \RegFile/_0253_ ;
wire \RegFile/_0254_ ;
wire \RegFile/_0255_ ;
wire \RegFile/_0256_ ;
wire \RegFile/_0257_ ;
wire \RegFile/_0258_ ;
wire \RegFile/_0259_ ;
wire \RegFile/_0260_ ;
wire \RegFile/_0261_ ;
wire \RegFile/_0262_ ;
wire \RegFile/_0263_ ;
wire \RegFile/_0264_ ;
wire \RegFile/_0265_ ;
wire \RegFile/_0266_ ;
wire \RegFile/_0267_ ;
wire \RegFile/_0268_ ;
wire \RegFile/_0269_ ;
wire \RegFile/_0270_ ;
wire \RegFile/_0271_ ;
wire \RegFile/_0272_ ;
wire \RegFile/_0273_ ;
wire \RegFile/_0274_ ;
wire \RegFile/_0275_ ;
wire \RegFile/_0276_ ;
wire \RegFile/_0277_ ;
wire \RegFile/_0278_ ;
wire \RegFile/_0279_ ;
wire \RegFile/_0280_ ;
wire \RegFile/_0281_ ;
wire \RegFile/_0282_ ;
wire \RegFile/_0283_ ;
wire \RegFile/_0284_ ;
wire \RegFile/_0285_ ;
wire \RegFile/_0286_ ;
wire \RegFile/_0287_ ;
wire \RegFile/_0288_ ;
wire \RegFile/_0289_ ;
wire \RegFile/_0290_ ;
wire \RegFile/_0291_ ;
wire \RegFile/_0292_ ;
wire \RegFile/_0293_ ;
wire \RegFile/_0294_ ;
wire \RegFile/_0295_ ;
wire \RegFile/_0296_ ;
wire \RegFile/_0297_ ;
wire \RegFile/_0298_ ;
wire \RegFile/_0299_ ;
wire \RegFile/_0300_ ;
wire \RegFile/_0301_ ;
wire \RegFile/_0302_ ;
wire \RegFile/_0303_ ;
wire \RegFile/_0304_ ;
wire \RegFile/_0305_ ;
wire \RegFile/_0306_ ;
wire \RegFile/_0307_ ;
wire \RegFile/_0308_ ;
wire \RegFile/_0309_ ;
wire \RegFile/_0310_ ;
wire \RegFile/_0311_ ;
wire \RegFile/_0312_ ;
wire \RegFile/_0313_ ;
wire \RegFile/_0314_ ;
wire \RegFile/_0315_ ;
wire \RegFile/_0316_ ;
wire \RegFile/_0317_ ;
wire \RegFile/_0318_ ;
wire \RegFile/_0319_ ;
wire \RegFile/_0320_ ;
wire \RegFile/_0321_ ;
wire \RegFile/_0322_ ;
wire \RegFile/_0323_ ;
wire \RegFile/_0324_ ;
wire \RegFile/_0325_ ;
wire \RegFile/_0326_ ;
wire \RegFile/_0327_ ;
wire \RegFile/_0328_ ;
wire \RegFile/_0329_ ;
wire \RegFile/_0330_ ;
wire \RegFile/_0331_ ;
wire \RegFile/_0332_ ;
wire \RegFile/_0333_ ;
wire \RegFile/_0334_ ;
wire \RegFile/_0335_ ;
wire \RegFile/_0336_ ;
wire \RegFile/_0337_ ;
wire \RegFile/_0338_ ;
wire \RegFile/_0339_ ;
wire \RegFile/_0340_ ;
wire \RegFile/_0341_ ;
wire \RegFile/_0342_ ;
wire \RegFile/_0343_ ;
wire \RegFile/_0344_ ;
wire \RegFile/_0345_ ;
wire \RegFile/_0346_ ;
wire \RegFile/_0347_ ;
wire \RegFile/_0348_ ;
wire \RegFile/_0349_ ;
wire \RegFile/_0350_ ;
wire \RegFile/_0351_ ;
wire \RegFile/_0352_ ;
wire \RegFile/_0353_ ;
wire \RegFile/_0354_ ;
wire \RegFile/_0355_ ;
wire \RegFile/_0356_ ;
wire \RegFile/_0357_ ;
wire \RegFile/_0358_ ;
wire \RegFile/_0359_ ;
wire \RegFile/_0360_ ;
wire \RegFile/_0361_ ;
wire \RegFile/_0362_ ;
wire \RegFile/_0363_ ;
wire \RegFile/_0364_ ;
wire \RegFile/_0365_ ;
wire \RegFile/_0366_ ;
wire \RegFile/_0367_ ;
wire \RegFile/_0368_ ;
wire \RegFile/_0369_ ;
wire \RegFile/_0370_ ;
wire \RegFile/_0371_ ;
wire \RegFile/_0372_ ;
wire \RegFile/_0373_ ;
wire \RegFile/_0374_ ;
wire \RegFile/_0375_ ;
wire \RegFile/_0376_ ;
wire \RegFile/_0377_ ;
wire \RegFile/_0378_ ;
wire \RegFile/_0379_ ;
wire \RegFile/_0380_ ;
wire \RegFile/_0381_ ;
wire \RegFile/_0382_ ;
wire \RegFile/_0383_ ;
wire \RegFile/_0384_ ;
wire \RegFile/_0385_ ;
wire \RegFile/_0386_ ;
wire \RegFile/_0387_ ;
wire \RegFile/_0388_ ;
wire \RegFile/_0389_ ;
wire \RegFile/_0390_ ;
wire \RegFile/_0391_ ;
wire \RegFile/_0392_ ;
wire \RegFile/_0393_ ;
wire \RegFile/_0394_ ;
wire \RegFile/_0395_ ;
wire \RegFile/_0396_ ;
wire \RegFile/_0397_ ;
wire \RegFile/_0398_ ;
wire \RegFile/_0399_ ;
wire \RegFile/_0400_ ;
wire \RegFile/_0401_ ;
wire \RegFile/_0402_ ;
wire \RegFile/_0403_ ;
wire \RegFile/_0404_ ;
wire \RegFile/_0405_ ;
wire \RegFile/_0406_ ;
wire \RegFile/_0407_ ;
wire \RegFile/_0408_ ;
wire \RegFile/_0409_ ;
wire \RegFile/_0410_ ;
wire \RegFile/_0411_ ;
wire \RegFile/_0412_ ;
wire \RegFile/_0413_ ;
wire \RegFile/_0414_ ;
wire \RegFile/_0415_ ;
wire \RegFile/_0416_ ;
wire \RegFile/_0417_ ;
wire \RegFile/_0418_ ;
wire \RegFile/_0419_ ;
wire \RegFile/_0420_ ;
wire \RegFile/_0421_ ;
wire \RegFile/_0422_ ;
wire \RegFile/_0423_ ;
wire \RegFile/_0424_ ;
wire \RegFile/_0425_ ;
wire \RegFile/_0426_ ;
wire \RegFile/_0427_ ;
wire \RegFile/_0428_ ;
wire \RegFile/_0429_ ;
wire \RegFile/_0430_ ;
wire \RegFile/_0431_ ;
wire \RegFile/_0432_ ;
wire \RegFile/_0433_ ;
wire \RegFile/_0434_ ;
wire \RegFile/_0435_ ;
wire \RegFile/_0436_ ;
wire \RegFile/_0437_ ;
wire \RegFile/_0438_ ;
wire \RegFile/_0439_ ;
wire \RegFile/_0440_ ;
wire \RegFile/_0441_ ;
wire \RegFile/_0442_ ;
wire \RegFile/_0443_ ;
wire \RegFile/_0444_ ;
wire \RegFile/_0445_ ;
wire \RegFile/_0446_ ;
wire \RegFile/_0447_ ;
wire \RegFile/_0448_ ;
wire \RegFile/_0449_ ;
wire \RegFile/_0450_ ;
wire \RegFile/_0451_ ;
wire \RegFile/_0452_ ;
wire \RegFile/_0453_ ;
wire \RegFile/_0454_ ;
wire \RegFile/_0455_ ;
wire \RegFile/_0456_ ;
wire \RegFile/_0457_ ;
wire \RegFile/_0458_ ;
wire \RegFile/_0459_ ;
wire \RegFile/_0460_ ;
wire \RegFile/_0461_ ;
wire \RegFile/_0462_ ;
wire \RegFile/_0463_ ;
wire \RegFile/_0464_ ;
wire \RegFile/_0465_ ;
wire \RegFile/_0466_ ;
wire \RegFile/_0467_ ;
wire \RegFile/_0468_ ;
wire \RegFile/_0469_ ;
wire \RegFile/_0470_ ;
wire \RegFile/_0471_ ;
wire \RegFile/_0472_ ;
wire \RegFile/_0473_ ;
wire \RegFile/_0474_ ;
wire \RegFile/_0475_ ;
wire \RegFile/_0476_ ;
wire \RegFile/_0477_ ;
wire \RegFile/_0478_ ;
wire \RegFile/_0479_ ;
wire \RegFile/_0480_ ;
wire \RegFile/_0481_ ;
wire \RegFile/_0482_ ;
wire \RegFile/_0483_ ;
wire \RegFile/_0484_ ;
wire \RegFile/_0485_ ;
wire \RegFile/_0486_ ;
wire \RegFile/_0487_ ;
wire \RegFile/_0488_ ;
wire \RegFile/_0489_ ;
wire \RegFile/_0490_ ;
wire \RegFile/_0491_ ;
wire \RegFile/_0492_ ;
wire \RegFile/_0493_ ;
wire \RegFile/_0494_ ;
wire \RegFile/_0495_ ;
wire \RegFile/_0496_ ;
wire \RegFile/_0497_ ;
wire \RegFile/_0498_ ;
wire \RegFile/_0499_ ;
wire \RegFile/_0500_ ;
wire \RegFile/_0501_ ;
wire \RegFile/_0502_ ;
wire \RegFile/_0503_ ;
wire \RegFile/_0504_ ;
wire \RegFile/_0505_ ;
wire \RegFile/_0506_ ;
wire \RegFile/_0507_ ;
wire \RegFile/_0508_ ;
wire \RegFile/_0509_ ;
wire \RegFile/_0510_ ;
wire \RegFile/_0511_ ;
wire \RegFile/_0512_ ;
wire \RegFile/_0513_ ;
wire \RegFile/_0514_ ;
wire \RegFile/_0515_ ;
wire \RegFile/_0516_ ;
wire \RegFile/_0517_ ;
wire \RegFile/_0518_ ;
wire \RegFile/_0519_ ;
wire \RegFile/_0520_ ;
wire \RegFile/_0521_ ;
wire \RegFile/_0522_ ;
wire \RegFile/_0523_ ;
wire \RegFile/_0524_ ;
wire \RegFile/_0525_ ;
wire \RegFile/_0526_ ;
wire \RegFile/_0527_ ;
wire \RegFile/_0528_ ;
wire \RegFile/_0529_ ;
wire \RegFile/_0530_ ;
wire \RegFile/_0531_ ;
wire \RegFile/_0532_ ;
wire \RegFile/_0533_ ;
wire \RegFile/_0534_ ;
wire \RegFile/_0535_ ;
wire \RegFile/_0536_ ;
wire \RegFile/_0537_ ;
wire \RegFile/_0538_ ;
wire \RegFile/_0539_ ;
wire \RegFile/_0540_ ;
wire \RegFile/_0541_ ;
wire \RegFile/_0542_ ;
wire \RegFile/_0543_ ;
wire \RegFile/_0544_ ;
wire \RegFile/_0545_ ;
wire \RegFile/_0546_ ;
wire \RegFile/_0547_ ;
wire \RegFile/_0548_ ;
wire \RegFile/_0549_ ;
wire \RegFile/_0550_ ;
wire \RegFile/_0551_ ;
wire \RegFile/_0552_ ;
wire \RegFile/_0553_ ;
wire \RegFile/_0554_ ;
wire \RegFile/_0555_ ;
wire \RegFile/_0556_ ;
wire \RegFile/_0557_ ;
wire \RegFile/_0558_ ;
wire \RegFile/_0559_ ;
wire \RegFile/_0560_ ;
wire \RegFile/_0561_ ;
wire \RegFile/_0562_ ;
wire \RegFile/_0563_ ;
wire \RegFile/_0564_ ;
wire \RegFile/_0565_ ;
wire \RegFile/_0566_ ;
wire \RegFile/_0567_ ;
wire \RegFile/_0568_ ;
wire \RegFile/_0569_ ;
wire \RegFile/_0570_ ;
wire \RegFile/_0571_ ;
wire \RegFile/_0572_ ;
wire \RegFile/_0573_ ;
wire \RegFile/_0574_ ;
wire \RegFile/_0575_ ;
wire \RegFile/_0576_ ;
wire \RegFile/_0577_ ;
wire \RegFile/_0578_ ;
wire \RegFile/_0579_ ;
wire \RegFile/_0580_ ;
wire \RegFile/_0581_ ;
wire \RegFile/_0582_ ;
wire \RegFile/_0583_ ;
wire \RegFile/_0584_ ;
wire \RegFile/_0585_ ;
wire \RegFile/_0586_ ;
wire \RegFile/_0587_ ;
wire \RegFile/_0588_ ;
wire \RegFile/_0589_ ;
wire \RegFile/_0590_ ;
wire \RegFile/_0591_ ;
wire \RegFile/_0592_ ;
wire \RegFile/_0593_ ;
wire \RegFile/_0594_ ;
wire \RegFile/_0595_ ;
wire \RegFile/_0596_ ;
wire \RegFile/_0597_ ;
wire \RegFile/_0598_ ;
wire \RegFile/_0599_ ;
wire \RegFile/_0600_ ;
wire \RegFile/_0601_ ;
wire \RegFile/_0602_ ;
wire \RegFile/_0603_ ;
wire \RegFile/_0604_ ;
wire \RegFile/_0605_ ;
wire \RegFile/_0606_ ;
wire \RegFile/_0607_ ;
wire \RegFile/_0608_ ;
wire \RegFile/_0609_ ;
wire \RegFile/_0610_ ;
wire \RegFile/_0611_ ;
wire \RegFile/_0612_ ;
wire \RegFile/_0613_ ;
wire \RegFile/_0614_ ;
wire \RegFile/_0615_ ;
wire \RegFile/_0616_ ;
wire \RegFile/_0617_ ;
wire \RegFile/_0618_ ;
wire \RegFile/_0619_ ;
wire \RegFile/_0620_ ;
wire \RegFile/_0621_ ;
wire \RegFile/_0622_ ;
wire \RegFile/_0623_ ;
wire \RegFile/_0624_ ;
wire \RegFile/_0625_ ;
wire \RegFile/_0626_ ;
wire \RegFile/_0627_ ;
wire \RegFile/_0628_ ;
wire \RegFile/_0629_ ;
wire \RegFile/_0630_ ;
wire \RegFile/_0631_ ;
wire \RegFile/_0632_ ;
wire \RegFile/_0633_ ;
wire \RegFile/_0634_ ;
wire \RegFile/_0635_ ;
wire \RegFile/_0636_ ;
wire \RegFile/_0637_ ;
wire \RegFile/_0638_ ;
wire \RegFile/_0639_ ;
wire \RegFile/_0640_ ;
wire \RegFile/_0641_ ;
wire \RegFile/_0642_ ;
wire \RegFile/_0643_ ;
wire \RegFile/_0644_ ;
wire \RegFile/_0645_ ;
wire \RegFile/_0646_ ;
wire \RegFile/_0647_ ;
wire \RegFile/_0648_ ;
wire \RegFile/_0649_ ;
wire \RegFile/_0650_ ;
wire \RegFile/_0651_ ;
wire \RegFile/_0652_ ;
wire \RegFile/_0653_ ;
wire \RegFile/_0654_ ;
wire \RegFile/_0655_ ;
wire \RegFile/_0656_ ;
wire \RegFile/_0657_ ;
wire \RegFile/_0658_ ;
wire \RegFile/_0659_ ;
wire \RegFile/_0660_ ;
wire \RegFile/_0661_ ;
wire \RegFile/_0662_ ;
wire \RegFile/_0663_ ;
wire \RegFile/_0664_ ;
wire \RegFile/_0665_ ;
wire \RegFile/_0666_ ;
wire \RegFile/_0667_ ;
wire \RegFile/_0668_ ;
wire \RegFile/_0669_ ;
wire \RegFile/_0670_ ;
wire \RegFile/_0671_ ;
wire \RegFile/_0672_ ;
wire \RegFile/_0673_ ;
wire \RegFile/_0674_ ;
wire \RegFile/_0675_ ;
wire \RegFile/_0676_ ;
wire \RegFile/_0677_ ;
wire \RegFile/_0678_ ;
wire \RegFile/_0679_ ;
wire \RegFile/_0680_ ;
wire \RegFile/_0681_ ;
wire \RegFile/_0682_ ;
wire \RegFile/_0683_ ;
wire \RegFile/_0684_ ;
wire \RegFile/_0685_ ;
wire \RegFile/_0686_ ;
wire \RegFile/_0687_ ;
wire \RegFile/_0688_ ;
wire \RegFile/_0689_ ;
wire \RegFile/_0690_ ;
wire \RegFile/_0691_ ;
wire \RegFile/_0692_ ;
wire \RegFile/_0693_ ;
wire \RegFile/_0694_ ;
wire \RegFile/_0695_ ;
wire \RegFile/_0696_ ;
wire \RegFile/_0697_ ;
wire \RegFile/_0698_ ;
wire \RegFile/_0699_ ;
wire \RegFile/_0700_ ;
wire \RegFile/_0701_ ;
wire \RegFile/_0702_ ;
wire \RegFile/_0703_ ;
wire \RegFile/_0704_ ;
wire \RegFile/_0705_ ;
wire \RegFile/_0706_ ;
wire \RegFile/_0707_ ;
wire \RegFile/_0708_ ;
wire \RegFile/_0709_ ;
wire \RegFile/_0710_ ;
wire \RegFile/_0711_ ;
wire \RegFile/_0712_ ;
wire \RegFile/_0713_ ;
wire \RegFile/_0714_ ;
wire \RegFile/_0715_ ;
wire \RegFile/_0716_ ;
wire \RegFile/_0717_ ;
wire \RegFile/_0718_ ;
wire \RegFile/_0719_ ;
wire \RegFile/_0720_ ;
wire \RegFile/_0721_ ;
wire \RegFile/_0722_ ;
wire \RegFile/_0723_ ;
wire \RegFile/_0724_ ;
wire \RegFile/_0725_ ;
wire \RegFile/_0726_ ;
wire \RegFile/_0727_ ;
wire \RegFile/_0728_ ;
wire \RegFile/_0729_ ;
wire \RegFile/_0730_ ;
wire \RegFile/_0731_ ;
wire \RegFile/_0732_ ;
wire \RegFile/_0733_ ;
wire \RegFile/_0734_ ;
wire \RegFile/_0735_ ;
wire \RegFile/_0736_ ;
wire \RegFile/_0737_ ;
wire \RegFile/_0738_ ;
wire \RegFile/_0739_ ;
wire \RegFile/_0740_ ;
wire \RegFile/_0741_ ;
wire \RegFile/_0742_ ;
wire \RegFile/_0743_ ;
wire \RegFile/_0744_ ;
wire \RegFile/_0745_ ;
wire \RegFile/_0746_ ;
wire \RegFile/_0747_ ;
wire \RegFile/_0748_ ;
wire \RegFile/_0749_ ;
wire \RegFile/_0750_ ;
wire \RegFile/_0751_ ;
wire \RegFile/_0752_ ;
wire \RegFile/_0753_ ;
wire \RegFile/_0754_ ;
wire \RegFile/_0755_ ;
wire \RegFile/_0756_ ;
wire \RegFile/_0757_ ;
wire \RegFile/_0758_ ;
wire \RegFile/_0759_ ;
wire \RegFile/_0760_ ;
wire \RegFile/_0761_ ;
wire \RegFile/_0762_ ;
wire \RegFile/_0763_ ;
wire \RegFile/_0764_ ;
wire \RegFile/_0765_ ;
wire \RegFile/_0766_ ;
wire \RegFile/_0767_ ;
wire \RegFile/_0768_ ;
wire \RegFile/_0769_ ;
wire \RegFile/_0770_ ;
wire \RegFile/_0771_ ;
wire \RegFile/_0772_ ;
wire \RegFile/_0773_ ;
wire \RegFile/_0774_ ;
wire \RegFile/_0775_ ;
wire \RegFile/_0776_ ;
wire \RegFile/_0777_ ;
wire \RegFile/_0778_ ;
wire \RegFile/_0779_ ;
wire \RegFile/_0780_ ;
wire \RegFile/_0781_ ;
wire \RegFile/_0782_ ;
wire \RegFile/_0783_ ;
wire \RegFile/_0784_ ;
wire \RegFile/_0785_ ;
wire \RegFile/_0786_ ;
wire \RegFile/_0787_ ;
wire \RegFile/_0788_ ;
wire \RegFile/_0789_ ;
wire \RegFile/_0790_ ;
wire \RegFile/_0791_ ;
wire \RegFile/_0792_ ;
wire \RegFile/_0793_ ;
wire \RegFile/_0794_ ;
wire \RegFile/_0795_ ;
wire \RegFile/_0796_ ;
wire \RegFile/_0797_ ;
wire \RegFile/_0798_ ;
wire \RegFile/_0799_ ;
wire \RegFile/_0800_ ;
wire \RegFile/_0801_ ;
wire \RegFile/_0802_ ;
wire \RegFile/_0803_ ;
wire \RegFile/_0804_ ;
wire \RegFile/_0805_ ;
wire \RegFile/_0806_ ;
wire \RegFile/_0807_ ;
wire \RegFile/_0808_ ;
wire \RegFile/_0809_ ;
wire \RegFile/_0810_ ;
wire \RegFile/_0811_ ;
wire \RegFile/_0812_ ;
wire \RegFile/_0813_ ;
wire \RegFile/_0814_ ;
wire \RegFile/_0815_ ;
wire \RegFile/_0816_ ;
wire \RegFile/_0817_ ;
wire \RegFile/_0818_ ;
wire \RegFile/_0819_ ;
wire \RegFile/_0820_ ;
wire \RegFile/_0821_ ;
wire \RegFile/_0822_ ;
wire \RegFile/_0823_ ;
wire \RegFile/_0824_ ;
wire \RegFile/_0825_ ;
wire \RegFile/_0826_ ;
wire \RegFile/_0827_ ;
wire \RegFile/_0828_ ;
wire \RegFile/_0829_ ;
wire \RegFile/_0830_ ;
wire \RegFile/_0831_ ;
wire \RegFile/_0832_ ;
wire \RegFile/_0833_ ;
wire \RegFile/_0834_ ;
wire \RegFile/_0835_ ;
wire \RegFile/_0836_ ;
wire \RegFile/_0837_ ;
wire \RegFile/_0838_ ;
wire \RegFile/_0839_ ;
wire \RegFile/_0840_ ;
wire \RegFile/_0841_ ;
wire \RegFile/_0842_ ;
wire \RegFile/_0843_ ;
wire \RegFile/_0844_ ;
wire \RegFile/_0845_ ;
wire \RegFile/_0846_ ;
wire \RegFile/_0847_ ;
wire \RegFile/_0848_ ;
wire \RegFile/_0849_ ;
wire \RegFile/_0850_ ;
wire \RegFile/_0851_ ;
wire \RegFile/_0852_ ;
wire \RegFile/_0853_ ;
wire \RegFile/_0854_ ;
wire \RegFile/_0855_ ;
wire \RegFile/_0856_ ;
wire \RegFile/_0857_ ;
wire \RegFile/_0858_ ;
wire \RegFile/_0859_ ;
wire \RegFile/_0860_ ;
wire \RegFile/_0861_ ;
wire \RegFile/_0862_ ;
wire \RegFile/_0863_ ;
wire \RegFile/_0864_ ;
wire \RegFile/_0865_ ;
wire \RegFile/_0866_ ;
wire \RegFile/_0867_ ;
wire \RegFile/_0868_ ;
wire \RegFile/_0869_ ;
wire \RegFile/_0870_ ;
wire \RegFile/_0871_ ;
wire \RegFile/_0872_ ;
wire \RegFile/_0873_ ;
wire \RegFile/_0874_ ;
wire \RegFile/_0875_ ;
wire \RegFile/_0876_ ;
wire \RegFile/_0877_ ;
wire \RegFile/_0878_ ;
wire \RegFile/_0879_ ;
wire \RegFile/_0880_ ;
wire \RegFile/_0881_ ;
wire \RegFile/_0882_ ;
wire \RegFile/_0883_ ;
wire \RegFile/_0884_ ;
wire \RegFile/_0885_ ;
wire \RegFile/_0886_ ;
wire \RegFile/_0887_ ;
wire \RegFile/_0888_ ;
wire \RegFile/_0889_ ;
wire \RegFile/_0890_ ;
wire \RegFile/_0891_ ;
wire \RegFile/_0892_ ;
wire \RegFile/_0893_ ;
wire \RegFile/_0894_ ;
wire \RegFile/_0895_ ;
wire \RegFile/_0896_ ;
wire \RegFile/_0897_ ;
wire \RegFile/_0898_ ;
wire \RegFile/_0899_ ;
wire \RegFile/_0900_ ;
wire \RegFile/_0901_ ;
wire \RegFile/_0902_ ;
wire \RegFile/_0903_ ;
wire \RegFile/_0904_ ;
wire \RegFile/_0905_ ;
wire \RegFile/_0906_ ;
wire \RegFile/_0907_ ;
wire \RegFile/_0908_ ;
wire \RegFile/_0909_ ;
wire \RegFile/_0910_ ;
wire \RegFile/_0911_ ;
wire \RegFile/_0912_ ;
wire \RegFile/_0913_ ;
wire \RegFile/_0914_ ;
wire \RegFile/_0915_ ;
wire \RegFile/_0916_ ;
wire \RegFile/_0917_ ;
wire \RegFile/_0918_ ;
wire \RegFile/_0919_ ;
wire \RegFile/_0920_ ;
wire \RegFile/_0921_ ;
wire \RegFile/_0922_ ;
wire \RegFile/_0923_ ;
wire \RegFile/_0924_ ;
wire \RegFile/_0925_ ;
wire \RegFile/_0926_ ;
wire \RegFile/_0927_ ;
wire \RegFile/_0928_ ;
wire \RegFile/_0929_ ;
wire \RegFile/_0930_ ;
wire \RegFile/_0931_ ;
wire \RegFile/_0932_ ;
wire \RegFile/_0933_ ;
wire \RegFile/_0934_ ;
wire \RegFile/_0935_ ;
wire \RegFile/_0936_ ;
wire \RegFile/_0937_ ;
wire \RegFile/_0938_ ;
wire \RegFile/_0939_ ;
wire \RegFile/_0940_ ;
wire \RegFile/_0941_ ;
wire \RegFile/_0942_ ;
wire \RegFile/_0943_ ;
wire \RegFile/_0944_ ;
wire \RegFile/_0945_ ;
wire \RegFile/_0946_ ;
wire \RegFile/_0947_ ;
wire \RegFile/_0948_ ;
wire \RegFile/_0949_ ;
wire \RegFile/_0950_ ;
wire \RegFile/_0951_ ;
wire \RegFile/_0952_ ;
wire \RegFile/_0953_ ;
wire \RegFile/_0954_ ;
wire \RegFile/_0955_ ;
wire \RegFile/_0956_ ;
wire \RegFile/_0957_ ;
wire \RegFile/_0958_ ;
wire \RegFile/_0959_ ;
wire \RegFile/_0960_ ;
wire \RegFile/_0961_ ;
wire \RegFile/_0962_ ;
wire \RegFile/_0963_ ;
wire \RegFile/_0964_ ;
wire \RegFile/_0965_ ;
wire \RegFile/_0966_ ;
wire \RegFile/_0967_ ;
wire \RegFile/_0968_ ;
wire \RegFile/_0969_ ;
wire \RegFile/_0970_ ;
wire \RegFile/_0971_ ;
wire \RegFile/_0972_ ;
wire \RegFile/_0973_ ;
wire \RegFile/_0974_ ;
wire \RegFile/_0975_ ;
wire \RegFile/_0976_ ;
wire \RegFile/_0977_ ;
wire \RegFile/_0978_ ;
wire \RegFile/_0979_ ;
wire \RegFile/_0980_ ;
wire \RegFile/_0981_ ;
wire \RegFile/_0982_ ;
wire \RegFile/_0983_ ;
wire \RegFile/_0984_ ;
wire \RegFile/_0985_ ;
wire \RegFile/_0986_ ;
wire \RegFile/_0987_ ;
wire \RegFile/_0988_ ;
wire \RegFile/_0989_ ;
wire \RegFile/_0990_ ;
wire \RegFile/_0991_ ;
wire \RegFile/_0992_ ;
wire \RegFile/_0993_ ;
wire \RegFile/_0994_ ;
wire \RegFile/_0995_ ;
wire \RegFile/_0996_ ;
wire \RegFile/_0997_ ;
wire \RegFile/_0998_ ;
wire \RegFile/_0999_ ;
wire \RegFile/_1000_ ;
wire \RegFile/_1001_ ;
wire \RegFile/_1002_ ;
wire \RegFile/_1003_ ;
wire \RegFile/_1004_ ;
wire \RegFile/_1005_ ;
wire \RegFile/_1006_ ;
wire \RegFile/_1007_ ;
wire \RegFile/_1008_ ;
wire \RegFile/_1009_ ;
wire \RegFile/_1010_ ;
wire \RegFile/_1011_ ;
wire \RegFile/_1012_ ;
wire \RegFile/_1013_ ;
wire \RegFile/_1014_ ;
wire \RegFile/_1015_ ;
wire \RegFile/_1016_ ;
wire \RegFile/_1017_ ;
wire \RegFile/_1018_ ;
wire \RegFile/_1019_ ;
wire \RegFile/_1020_ ;
wire \RegFile/_1021_ ;
wire \RegFile/_1022_ ;
wire \RegFile/_1023_ ;
wire \RegFile/_1024_ ;
wire \RegFile/_1025_ ;
wire \RegFile/_1026_ ;
wire \RegFile/_1027_ ;
wire \RegFile/_1028_ ;
wire \RegFile/_1029_ ;
wire \RegFile/_1030_ ;
wire \RegFile/_1031_ ;
wire \RegFile/_1032_ ;
wire \RegFile/_1033_ ;
wire \RegFile/_1034_ ;
wire \RegFile/_1035_ ;
wire \RegFile/_1036_ ;
wire \RegFile/_1037_ ;
wire \RegFile/_1038_ ;
wire \RegFile/_1039_ ;
wire \RegFile/_1040_ ;
wire \RegFile/_1041_ ;
wire \RegFile/_1042_ ;
wire \RegFile/_1043_ ;
wire \RegFile/_1044_ ;
wire \RegFile/_1045_ ;
wire \RegFile/_1046_ ;
wire \RegFile/_1047_ ;
wire \RegFile/_1048_ ;
wire \RegFile/_1049_ ;
wire \RegFile/_1050_ ;
wire \RegFile/_1051_ ;
wire \RegFile/_1052_ ;
wire \RegFile/_1053_ ;
wire \RegFile/_1054_ ;
wire \RegFile/_1055_ ;
wire \RegFile/_1056_ ;
wire \RegFile/_1057_ ;
wire \RegFile/_1058_ ;
wire \RegFile/_1059_ ;
wire \RegFile/_1060_ ;
wire \RegFile/_1061_ ;
wire \RegFile/_1062_ ;
wire \RegFile/_1063_ ;
wire \RegFile/_1064_ ;
wire \RegFile/_1065_ ;
wire \RegFile/_1066_ ;
wire \RegFile/_1067_ ;
wire \RegFile/_1068_ ;
wire \RegFile/_1069_ ;
wire \RegFile/_1070_ ;
wire \RegFile/_1071_ ;
wire \RegFile/_1072_ ;
wire \RegFile/_1073_ ;
wire \RegFile/_1074_ ;
wire \RegFile/_1075_ ;
wire \RegFile/_1076_ ;
wire \RegFile/_1077_ ;
wire \RegFile/_1078_ ;
wire \RegFile/_1079_ ;
wire \RegFile/_1080_ ;
wire \RegFile/_1081_ ;
wire \RegFile/_1082_ ;
wire \RegFile/_1083_ ;
wire \RegFile/_1084_ ;
wire \RegFile/_1085_ ;
wire \RegFile/_1086_ ;
wire \RegFile/_1087_ ;
wire \RegFile/_1088_ ;
wire \RegFile/_1089_ ;
wire \RegFile/_1090_ ;
wire \RegFile/_1091_ ;
wire \RegFile/_1092_ ;
wire \RegFile/_1093_ ;
wire \RegFile/_1094_ ;
wire \RegFile/_1095_ ;
wire \RegFile/_1096_ ;
wire \RegFile/_1097_ ;
wire \RegFile/_1098_ ;
wire \RegFile/_1099_ ;
wire \RegFile/_1100_ ;
wire \RegFile/_1101_ ;
wire \RegFile/_1102_ ;
wire \RegFile/_1103_ ;
wire \RegFile/_1104_ ;
wire \RegFile/_1105_ ;
wire \RegFile/_1106_ ;
wire \RegFile/_1107_ ;
wire \RegFile/_1108_ ;
wire \RegFile/_1109_ ;
wire \RegFile/_1110_ ;
wire \RegFile/_1111_ ;
wire \RegFile/_1112_ ;
wire \RegFile/_1113_ ;
wire \RegFile/_1114_ ;
wire \RegFile/_1115_ ;
wire \RegFile/_1116_ ;
wire \RegFile/_1117_ ;
wire \RegFile/_1118_ ;
wire \RegFile/_1119_ ;
wire \RegFile/_1120_ ;
wire \RegFile/_1121_ ;
wire \RegFile/_1122_ ;
wire \RegFile/_1123_ ;
wire \RegFile/_1124_ ;
wire \RegFile/_1125_ ;
wire \RegFile/_1126_ ;
wire \RegFile/_1127_ ;
wire \RegFile/_1128_ ;
wire \RegFile/_1129_ ;
wire \RegFile/_1130_ ;
wire \RegFile/_1131_ ;
wire \RegFile/_1132_ ;
wire \RegFile/_1133_ ;
wire \RegFile/_1134_ ;
wire \RegFile/_1135_ ;
wire \RegFile/_1136_ ;
wire \RegFile/_1137_ ;
wire \RegFile/_1138_ ;
wire \RegFile/_1139_ ;
wire \RegFile/_1140_ ;
wire \RegFile/_1141_ ;
wire \RegFile/_1142_ ;
wire \RegFile/_1143_ ;
wire \RegFile/_1144_ ;
wire \RegFile/_1145_ ;
wire \RegFile/_1146_ ;
wire \RegFile/_1147_ ;
wire \RegFile/_1148_ ;
wire \RegFile/_1149_ ;
wire \RegFile/_1150_ ;
wire \RegFile/_1151_ ;
wire \RegFile/_1152_ ;
wire \RegFile/_1153_ ;
wire \RegFile/_1154_ ;
wire \RegFile/_1155_ ;
wire \RegFile/_1156_ ;
wire \RegFile/_1157_ ;
wire \RegFile/_1158_ ;
wire \RegFile/_1159_ ;
wire \RegFile/_1160_ ;
wire \RegFile/_1161_ ;
wire \RegFile/_1162_ ;
wire \RegFile/_1163_ ;
wire \RegFile/_1164_ ;
wire \RegFile/_1165_ ;
wire \RegFile/_1166_ ;
wire \RegFile/_1167_ ;
wire \RegFile/_1168_ ;
wire \RegFile/_1169_ ;
wire \RegFile/_1170_ ;
wire \RegFile/_1171_ ;
wire \RegFile/_1172_ ;
wire \RegFile/_1173_ ;
wire \RegFile/_1174_ ;
wire \RegFile/_1175_ ;
wire \RegFile/_1176_ ;
wire \RegFile/_1177_ ;
wire \RegFile/_1178_ ;
wire \RegFile/_1179_ ;
wire \RegFile/_1180_ ;
wire \RegFile/_1181_ ;
wire \RegFile/_1182_ ;
wire \RegFile/_1183_ ;
wire \RegFile/_1184_ ;
wire \RegFile/_1185_ ;
wire \RegFile/_1186_ ;
wire \RegFile/_1187_ ;
wire \RegFile/_1188_ ;
wire \RegFile/_1189_ ;
wire \RegFile/_1190_ ;
wire \RegFile/_1191_ ;
wire \RegFile/_1192_ ;
wire \RegFile/_1193_ ;
wire \RegFile/_1194_ ;
wire \RegFile/_1195_ ;
wire \RegFile/_1196_ ;
wire \RegFile/_1197_ ;
wire \RegFile/_1198_ ;
wire \RegFile/_1199_ ;
wire \RegFile/_1200_ ;
wire \RegFile/_1201_ ;
wire \RegFile/_1202_ ;
wire \RegFile/_1203_ ;
wire \RegFile/_1204_ ;
wire \RegFile/_1205_ ;
wire \RegFile/_1206_ ;
wire \RegFile/_1207_ ;
wire \RegFile/_1208_ ;
wire \RegFile/_1209_ ;
wire \RegFile/_1210_ ;
wire \RegFile/_1211_ ;
wire \RegFile/_1212_ ;
wire \RegFile/_1213_ ;
wire \RegFile/_1214_ ;
wire \RegFile/_1215_ ;
wire \RegFile/_1216_ ;
wire \RegFile/_1217_ ;
wire \RegFile/_1218_ ;
wire \RegFile/_1219_ ;
wire \RegFile/_1220_ ;
wire \RegFile/_1221_ ;
wire \RegFile/_1222_ ;
wire \RegFile/_1223_ ;
wire \RegFile/_1224_ ;
wire \RegFile/_1225_ ;
wire \RegFile/_1226_ ;
wire \RegFile/_1227_ ;
wire \RegFile/_1228_ ;
wire \RegFile/_1229_ ;
wire \RegFile/_1230_ ;
wire \RegFile/_1231_ ;
wire \RegFile/_1232_ ;
wire \RegFile/_1233_ ;
wire \RegFile/_1234_ ;
wire \RegFile/_1235_ ;
wire \RegFile/_1236_ ;
wire \RegFile/_1237_ ;
wire \RegFile/_1238_ ;
wire \RegFile/_1239_ ;
wire \RegFile/_1240_ ;
wire \RegFile/_1241_ ;
wire \RegFile/_1242_ ;
wire \RegFile/_1243_ ;
wire \RegFile/_1244_ ;
wire \RegFile/_1245_ ;
wire \RegFile/_1246_ ;
wire \RegFile/_1247_ ;
wire \RegFile/_1248_ ;
wire \RegFile/_1249_ ;
wire \RegFile/_1250_ ;
wire \RegFile/_1251_ ;
wire \RegFile/_1252_ ;
wire \RegFile/_1253_ ;
wire \RegFile/_1254_ ;
wire \RegFile/_1255_ ;
wire \RegFile/_1256_ ;
wire \RegFile/_1257_ ;
wire \RegFile/_1258_ ;
wire \RegFile/_1259_ ;
wire \RegFile/_1260_ ;
wire \RegFile/_1261_ ;
wire \RegFile/_1262_ ;
wire \RegFile/_1263_ ;
wire \RegFile/_1264_ ;
wire \RegFile/_1265_ ;
wire \RegFile/_1266_ ;
wire \RegFile/_1267_ ;
wire \RegFile/_1268_ ;
wire \RegFile/_1269_ ;
wire \RegFile/_1270_ ;
wire \RegFile/_1271_ ;
wire \RegFile/_1272_ ;
wire \RegFile/_1273_ ;
wire \RegFile/_1274_ ;
wire \RegFile/_1275_ ;
wire \RegFile/_1276_ ;
wire \RegFile/_1277_ ;
wire \RegFile/_1278_ ;
wire \RegFile/_1279_ ;
wire \RegFile/_1280_ ;
wire \RegFile/_1281_ ;
wire \RegFile/_1282_ ;
wire \RegFile/_1283_ ;
wire \RegFile/_1284_ ;
wire \RegFile/_1285_ ;
wire \RegFile/_1286_ ;
wire \RegFile/_1287_ ;
wire \RegFile/_1288_ ;
wire \RegFile/_1289_ ;
wire \RegFile/_1290_ ;
wire \RegFile/_1291_ ;
wire \RegFile/_1292_ ;
wire \RegFile/_1293_ ;
wire \RegFile/_1294_ ;
wire \RegFile/_1295_ ;
wire \RegFile/_1296_ ;
wire \RegFile/_1297_ ;
wire \RegFile/_1298_ ;
wire \RegFile/_1299_ ;
wire \RegFile/_1300_ ;
wire \RegFile/_1301_ ;
wire \RegFile/_1302_ ;
wire \RegFile/_1303_ ;
wire \RegFile/_1304_ ;
wire \RegFile/_1305_ ;
wire \RegFile/_1306_ ;
wire \RegFile/_1307_ ;
wire \RegFile/_1308_ ;
wire \RegFile/_1309_ ;
wire \RegFile/_1310_ ;
wire \RegFile/_1311_ ;
wire \RegFile/_1312_ ;
wire \RegFile/_1313_ ;
wire \RegFile/_1314_ ;
wire \RegFile/_1315_ ;
wire \RegFile/_1316_ ;
wire \RegFile/_1317_ ;
wire \RegFile/_1318_ ;
wire \RegFile/_1319_ ;
wire \RegFile/_1320_ ;
wire \RegFile/_1321_ ;
wire \RegFile/_1322_ ;
wire \RegFile/_1323_ ;
wire \RegFile/_1324_ ;
wire \RegFile/_1325_ ;
wire \RegFile/_1326_ ;
wire \RegFile/_1327_ ;
wire \RegFile/_1328_ ;
wire \RegFile/_1329_ ;
wire \RegFile/_1330_ ;
wire \RegFile/_1331_ ;
wire \RegFile/_1332_ ;
wire \RegFile/_1333_ ;
wire \RegFile/_1334_ ;
wire \RegFile/_1335_ ;
wire \RegFile/_1336_ ;
wire \RegFile/_1337_ ;
wire \RegFile/_1338_ ;
wire \RegFile/_1339_ ;
wire \RegFile/_1340_ ;
wire \RegFile/_1341_ ;
wire \RegFile/_1342_ ;
wire \RegFile/_1343_ ;
wire \RegFile/_1344_ ;
wire \RegFile/_1345_ ;
wire \RegFile/_1346_ ;
wire \RegFile/_1347_ ;
wire \RegFile/_1348_ ;
wire \RegFile/_1349_ ;
wire \RegFile/_1350_ ;
wire \RegFile/_1351_ ;
wire \RegFile/_1352_ ;
wire \RegFile/_1353_ ;
wire \RegFile/_1354_ ;
wire \RegFile/_1355_ ;
wire \RegFile/_1356_ ;
wire \RegFile/_1357_ ;
wire \RegFile/_1358_ ;
wire \RegFile/_1359_ ;
wire \RegFile/_1360_ ;
wire \RegFile/_1361_ ;
wire \RegFile/_1362_ ;
wire \RegFile/_1363_ ;
wire \RegFile/_1364_ ;
wire \RegFile/_1365_ ;
wire \RegFile/_1366_ ;
wire \RegFile/_1367_ ;
wire \RegFile/_1368_ ;
wire \RegFile/_1369_ ;
wire \RegFile/_1370_ ;
wire \RegFile/_1371_ ;
wire \RegFile/_1372_ ;
wire \RegFile/_1373_ ;
wire \RegFile/_1374_ ;
wire \RegFile/_1375_ ;
wire \RegFile/_1376_ ;
wire \RegFile/_1377_ ;
wire \RegFile/_1378_ ;
wire \RegFile/_1379_ ;
wire \RegFile/_1380_ ;
wire \RegFile/_1381_ ;
wire \RegFile/_1382_ ;
wire \RegFile/_1383_ ;
wire \RegFile/_1384_ ;
wire \RegFile/_1385_ ;
wire \RegFile/_1386_ ;
wire \RegFile/_1387_ ;
wire \RegFile/_1388_ ;
wire \RegFile/_1389_ ;
wire \RegFile/_1390_ ;
wire \RegFile/_1391_ ;
wire \RegFile/_1392_ ;
wire \RegFile/_1393_ ;
wire \RegFile/_1394_ ;
wire \RegFile/_1395_ ;
wire \RegFile/_1396_ ;
wire \RegFile/_1397_ ;
wire \RegFile/_1398_ ;
wire \RegFile/_1399_ ;
wire \RegFile/_1400_ ;
wire \RegFile/_1401_ ;
wire \RegFile/_1402_ ;
wire \RegFile/_1403_ ;
wire \RegFile/_1404_ ;
wire \RegFile/_1405_ ;
wire \RegFile/_1406_ ;
wire \RegFile/_1407_ ;
wire \RegFile/_1408_ ;
wire \RegFile/_1409_ ;
wire \RegFile/_1410_ ;
wire \RegFile/_1411_ ;
wire \RegFile/_1412_ ;
wire \RegFile/_1413_ ;
wire \RegFile/_1414_ ;
wire \RegFile/_1415_ ;
wire \RegFile/_1416_ ;
wire \RegFile/_1417_ ;
wire \RegFile/_1418_ ;
wire \RegFile/_1419_ ;
wire \RegFile/_1420_ ;
wire \RegFile/_1421_ ;
wire \RegFile/_1422_ ;
wire \RegFile/_1423_ ;
wire \RegFile/_1424_ ;
wire \RegFile/_1425_ ;
wire \RegFile/_1426_ ;
wire \RegFile/_1427_ ;
wire \RegFile/_1428_ ;
wire \RegFile/_1429_ ;
wire \RegFile/_1430_ ;
wire \RegFile/_1431_ ;
wire \RegFile/_1432_ ;
wire \RegFile/_1433_ ;
wire \RegFile/_1434_ ;
wire \RegFile/_1435_ ;
wire \RegFile/_1436_ ;
wire \RegFile/_1437_ ;
wire \RegFile/_1438_ ;
wire \RegFile/_1439_ ;
wire \RegFile/_1440_ ;
wire \RegFile/_1441_ ;
wire \RegFile/_1442_ ;
wire \RegFile/_1443_ ;
wire \RegFile/_1444_ ;
wire \RegFile/_1445_ ;
wire \RegFile/_1446_ ;
wire \RegFile/_1447_ ;
wire \RegFile/_1448_ ;
wire \RegFile/_1449_ ;
wire \RegFile/_1450_ ;
wire \RegFile/_1451_ ;
wire \RegFile/_1452_ ;
wire \RegFile/_1453_ ;
wire \RegFile/_1454_ ;
wire \RegFile/_1455_ ;
wire \RegFile/_1456_ ;
wire \RegFile/_1457_ ;
wire \RegFile/_1458_ ;
wire \RegFile/_1459_ ;
wire \RegFile/_1460_ ;
wire \RegFile/_1461_ ;
wire \RegFile/_1462_ ;
wire \RegFile/_1463_ ;
wire \RegFile/_1464_ ;
wire \RegFile/_1465_ ;
wire \RegFile/_1466_ ;
wire \RegFile/_1467_ ;
wire \RegFile/_1468_ ;
wire \RegFile/_1469_ ;
wire \RegFile/_1470_ ;
wire \RegFile/_1471_ ;
wire \RegFile/_1472_ ;
wire \RegFile/_1473_ ;
wire \RegFile/_1474_ ;
wire \RegFile/_1475_ ;
wire \RegFile/_1476_ ;
wire \RegFile/_1477_ ;
wire \RegFile/_1478_ ;
wire \RegFile/_1479_ ;
wire \RegFile/_1480_ ;
wire \RegFile/_1481_ ;
wire \RegFile/_1482_ ;
wire \RegFile/_1483_ ;
wire \RegFile/_1484_ ;
wire \RegFile/_1485_ ;
wire \RegFile/_1486_ ;
wire \RegFile/_1487_ ;
wire \RegFile/_1488_ ;
wire \RegFile/_1489_ ;
wire \RegFile/_1490_ ;
wire \RegFile/_1491_ ;
wire \RegFile/_1492_ ;
wire \RegFile/_1493_ ;
wire \RegFile/_1494_ ;
wire \RegFile/_1495_ ;
wire \RegFile/_1496_ ;
wire \RegFile/_1497_ ;
wire \RegFile/_1498_ ;
wire \RegFile/_1499_ ;
wire \RegFile/_1500_ ;
wire \RegFile/_1501_ ;
wire \RegFile/_1502_ ;
wire \RegFile/_1503_ ;
wire \RegFile/_1504_ ;
wire \RegFile/_1505_ ;
wire \RegFile/_1506_ ;
wire \RegFile/_1507_ ;
wire \RegFile/_1508_ ;
wire \RegFile/_1509_ ;
wire \RegFile/_1510_ ;
wire \RegFile/_1511_ ;
wire \RegFile/_1512_ ;
wire \RegFile/_1513_ ;
wire \RegFile/_1514_ ;
wire \RegFile/_1515_ ;
wire \RegFile/_1516_ ;
wire \RegFile/_1517_ ;
wire \RegFile/_1518_ ;
wire \RegFile/_1519_ ;
wire \RegFile/_1520_ ;
wire \RegFile/_1521_ ;
wire \RegFile/_1522_ ;
wire \RegFile/_1523_ ;
wire \RegFile/_1524_ ;
wire \RegFile/_1525_ ;
wire \RegFile/_1526_ ;
wire \RegFile/_1527_ ;
wire \RegFile/_1528_ ;
wire \RegFile/_1529_ ;
wire \RegFile/_1530_ ;
wire \RegFile/_1531_ ;
wire \RegFile/_1532_ ;
wire \RegFile/_1533_ ;
wire \RegFile/_1534_ ;
wire \RegFile/_1535_ ;
wire \RegFile/_1536_ ;
wire \RegFile/_1537_ ;
wire \RegFile/_1538_ ;
wire \RegFile/_1539_ ;
wire \RegFile/_1540_ ;
wire \RegFile/_1541_ ;
wire \RegFile/_1542_ ;
wire \RegFile/_1543_ ;
wire \RegFile/_1544_ ;
wire \RegFile/_1545_ ;
wire \RegFile/_1546_ ;
wire \RegFile/_1547_ ;
wire \RegFile/_1548_ ;
wire \RegFile/_1549_ ;
wire \RegFile/_1550_ ;
wire \RegFile/_1551_ ;
wire \RegFile/_1552_ ;
wire \RegFile/_1553_ ;
wire \RegFile/_1554_ ;
wire \RegFile/_1555_ ;
wire \RegFile/_1556_ ;
wire \RegFile/_1557_ ;
wire \RegFile/_1558_ ;
wire \RegFile/_1559_ ;
wire \RegFile/_1560_ ;
wire \RegFile/_1561_ ;
wire \RegFile/_1562_ ;
wire \RegFile/_1563_ ;
wire \RegFile/_1564_ ;
wire \RegFile/_1565_ ;
wire \RegFile/_1566_ ;
wire \RegFile/_1567_ ;
wire \RegFile/_1568_ ;
wire \RegFile/_1569_ ;
wire \RegFile/_1570_ ;
wire \RegFile/_1571_ ;
wire \RegFile/_1572_ ;
wire \RegFile/_1573_ ;
wire \RegFile/_1574_ ;
wire \RegFile/_1575_ ;
wire \RegFile/_1576_ ;
wire \RegFile/_1577_ ;
wire \RegFile/_1578_ ;
wire \RegFile/_1579_ ;
wire \RegFile/_1580_ ;
wire \RegFile/_1581_ ;
wire \RegFile/_1582_ ;
wire \RegFile/_1583_ ;
wire \RegFile/_1584_ ;
wire \RegFile/_1585_ ;
wire \RegFile/_1586_ ;
wire \RegFile/_1587_ ;
wire \RegFile/_1588_ ;
wire \RegFile/_1589_ ;
wire \RegFile/_1590_ ;
wire \RegFile/_1591_ ;
wire \RegFile/_1592_ ;
wire \RegFile/_1593_ ;
wire \RegFile/_1594_ ;
wire \RegFile/_1595_ ;
wire \RegFile/_1596_ ;
wire \RegFile/_1597_ ;
wire \RegFile/_1598_ ;
wire \RegFile/_1599_ ;
wire \RegFile/_1600_ ;
wire \RegFile/_1601_ ;
wire \RegFile/_1602_ ;
wire \RegFile/_1603_ ;
wire \RegFile/_1604_ ;
wire \RegFile/_1605_ ;
wire \RegFile/_1606_ ;
wire \RegFile/_1607_ ;
wire \RegFile/_1608_ ;
wire \RegFile/_1609_ ;
wire \RegFile/_1610_ ;
wire \RegFile/_1611_ ;
wire \RegFile/_1612_ ;
wire \RegFile/_1613_ ;
wire \RegFile/_1614_ ;
wire \RegFile/_1615_ ;
wire \RegFile/_1616_ ;
wire \RegFile/_1617_ ;
wire \RegFile/_1618_ ;
wire \RegFile/_1619_ ;
wire \RegFile/_1620_ ;
wire \RegFile/_1621_ ;
wire \RegFile/_1622_ ;
wire \RegFile/_1623_ ;
wire \RegFile/_1624_ ;
wire \RegFile/_1625_ ;
wire \RegFile/_1626_ ;
wire \RegFile/_1627_ ;
wire \RegFile/_1628_ ;
wire \RegFile/_1629_ ;
wire \RegFile/_1630_ ;
wire \RegFile/_1631_ ;
wire \RegFile/_1632_ ;
wire \RegFile/_1633_ ;
wire \RegFile/_1634_ ;
wire \RegFile/_1635_ ;
wire \RegFile/_1636_ ;
wire \RegFile/_1637_ ;
wire \RegFile/_1638_ ;
wire \RegFile/_1639_ ;
wire \RegFile/_1640_ ;
wire \RegFile/_1641_ ;
wire \RegFile/_1642_ ;
wire \RegFile/_1643_ ;
wire \RegFile/_1644_ ;
wire \RegFile/_1645_ ;
wire \RegFile/_1646_ ;
wire \RegFile/_1647_ ;
wire \RegFile/_1648_ ;
wire \RegFile/_1649_ ;
wire \RegFile/_1650_ ;
wire \RegFile/_1651_ ;
wire \RegFile/_1652_ ;
wire \RegFile/_1653_ ;
wire \RegFile/_1654_ ;
wire \RegFile/_1655_ ;
wire \RegFile/_1656_ ;
wire \RegFile/_1657_ ;
wire \RegFile/_1658_ ;
wire \RegFile/_1659_ ;
wire \RegFile/_1660_ ;
wire \RegFile/_1661_ ;
wire \RegFile/_1662_ ;
wire \RegFile/_1663_ ;
wire \RegFile/_1664_ ;
wire \RegFile/_1665_ ;
wire \RegFile/_1666_ ;
wire \RegFile/_1667_ ;
wire \RegFile/_1668_ ;
wire \RegFile/_1669_ ;
wire \RegFile/_1670_ ;
wire \RegFile/_1671_ ;
wire \RegFile/_1672_ ;
wire \RegFile/_1673_ ;
wire \RegFile/_1674_ ;
wire \RegFile/_1675_ ;
wire \RegFile/_1676_ ;
wire \RegFile/_1677_ ;
wire \RegFile/_1678_ ;
wire \RegFile/_1679_ ;
wire \RegFile/_1680_ ;
wire \RegFile/_1681_ ;
wire \RegFile/_1682_ ;
wire \RegFile/_1683_ ;
wire \RegFile/_1684_ ;
wire \RegFile/_1685_ ;
wire \RegFile/_1686_ ;
wire \RegFile/_1687_ ;
wire \RegFile/_1688_ ;
wire \RegFile/_1689_ ;
wire \RegFile/_1690_ ;
wire \RegFile/_1691_ ;
wire \RegFile/_1692_ ;
wire \RegFile/_1693_ ;
wire \RegFile/_1694_ ;
wire \RegFile/_1695_ ;
wire \RegFile/_1696_ ;
wire \RegFile/_1697_ ;
wire \RegFile/_1698_ ;
wire \RegFile/_1699_ ;
wire \RegFile/_1700_ ;
wire \RegFile/_1701_ ;
wire \RegFile/_1702_ ;
wire \RegFile/_1703_ ;
wire \RegFile/_1704_ ;
wire \RegFile/_1705_ ;
wire \RegFile/_1706_ ;
wire \RegFile/_1707_ ;
wire \RegFile/_1708_ ;
wire \RegFile/_1709_ ;
wire \RegFile/_1710_ ;
wire \RegFile/_1711_ ;
wire \RegFile/_1712_ ;
wire \RegFile/_1713_ ;
wire \RegFile/_1714_ ;
wire \RegFile/_1715_ ;
wire \RegFile/_1716_ ;
wire \RegFile/_1717_ ;
wire \RegFile/_1718_ ;
wire \RegFile/_1719_ ;
wire \RegFile/_1720_ ;
wire \RegFile/_1721_ ;
wire \RegFile/_1722_ ;
wire \RegFile/_1723_ ;
wire \RegFile/_1724_ ;
wire \RegFile/_1725_ ;
wire \RegFile/_1726_ ;
wire \RegFile/_1727_ ;
wire \RegFile/_1728_ ;
wire \RegFile/_1729_ ;
wire \RegFile/_1730_ ;
wire \RegFile/_1731_ ;
wire \RegFile/_1732_ ;
wire \RegFile/_1733_ ;
wire \RegFile/_1734_ ;
wire \RegFile/_1735_ ;
wire \RegFile/_1736_ ;
wire \RegFile/_1737_ ;
wire \RegFile/_1738_ ;
wire \RegFile/_1739_ ;
wire \RegFile/_1740_ ;
wire \RegFile/_1741_ ;
wire \RegFile/_1742_ ;
wire \RegFile/_1743_ ;
wire \RegFile/_1744_ ;
wire \RegFile/_1745_ ;
wire \RegFile/_1746_ ;
wire \RegFile/_1747_ ;
wire \RegFile/_1748_ ;
wire \RegFile/_1749_ ;
wire \RegFile/_1750_ ;
wire \RegFile/_1751_ ;
wire \RegFile/_1752_ ;
wire \RegFile/_1753_ ;
wire \RegFile/_1754_ ;
wire \RegFile/_1755_ ;
wire \RegFile/_1756_ ;
wire \RegFile/_1757_ ;
wire \RegFile/_1758_ ;
wire \RegFile/_1759_ ;
wire \RegFile/_1760_ ;
wire \RegFile/_1761_ ;
wire \RegFile/_1762_ ;
wire \RegFile/_1763_ ;
wire \RegFile/_1764_ ;
wire \RegFile/_1765_ ;
wire \RegFile/_1766_ ;
wire \RegFile/_1767_ ;
wire \RegFile/_1768_ ;
wire \RegFile/_1769_ ;
wire \RegFile/_1770_ ;
wire \RegFile/_1771_ ;
wire \RegFile/_1772_ ;
wire \RegFile/_1773_ ;
wire \RegFile/_1774_ ;
wire \RegFile/_1775_ ;
wire \RegFile/_1776_ ;
wire \RegFile/_1777_ ;
wire \RegFile/_1778_ ;
wire \RegFile/_1779_ ;
wire \RegFile/_1780_ ;
wire \RegFile/_1781_ ;
wire \RegFile/_1782_ ;
wire \RegFile/_1783_ ;
wire \RegFile/_1784_ ;
wire \RegFile/_1785_ ;
wire \RegFile/_1786_ ;
wire \RegFile/_1787_ ;
wire \RegFile/_1788_ ;
wire \RegFile/_1789_ ;
wire \RegFile/_1790_ ;
wire \RegFile/_1791_ ;
wire \RegFile/_1792_ ;
wire \RegFile/_1793_ ;
wire \RegFile/_1794_ ;
wire \RegFile/_1795_ ;
wire \RegFile/_1796_ ;
wire \RegFile/_1797_ ;
wire \RegFile/_1798_ ;
wire \RegFile/_1799_ ;
wire \RegFile/_1800_ ;
wire \RegFile/_1801_ ;
wire \RegFile/_1802_ ;
wire \RegFile/_1803_ ;
wire \RegFile/_1804_ ;
wire \RegFile/_1805_ ;
wire \RegFile/_1806_ ;
wire \RegFile/_1807_ ;
wire \RegFile/_1808_ ;
wire \RegFile/_1809_ ;
wire \RegFile/_1810_ ;
wire \RegFile/_1811_ ;
wire \RegFile/_1812_ ;
wire \RegFile/_1813_ ;
wire \RegFile/_1814_ ;
wire \RegFile/_1815_ ;
wire \RegFile/_1816_ ;
wire \RegFile/_1817_ ;
wire \RegFile/_1818_ ;
wire \RegFile/_1819_ ;
wire \RegFile/_1820_ ;
wire \RegFile/_1821_ ;
wire \RegFile/_1822_ ;
wire \RegFile/_1823_ ;
wire \RegFile/_1824_ ;
wire \RegFile/_1825_ ;
wire \RegFile/_1826_ ;
wire \RegFile/_1827_ ;
wire \RegFile/_1828_ ;
wire \RegFile/_1829_ ;
wire \RegFile/_1830_ ;
wire \RegFile/_1831_ ;
wire \RegFile/_1832_ ;
wire \RegFile/_1833_ ;
wire \RegFile/_1834_ ;
wire \RegFile/_1835_ ;
wire \RegFile/_1836_ ;
wire \RegFile/_1837_ ;
wire \RegFile/_1838_ ;
wire \RegFile/_1839_ ;
wire \RegFile/_1840_ ;
wire \RegFile/_1841_ ;
wire \RegFile/_1842_ ;
wire \RegFile/_1843_ ;
wire \RegFile/_1844_ ;
wire \RegFile/_1845_ ;
wire \RegFile/_1846_ ;
wire \RegFile/_1847_ ;
wire \RegFile/_1848_ ;
wire \RegFile/_1849_ ;
wire \RegFile/_1850_ ;
wire \RegFile/_1851_ ;
wire \RegFile/_1852_ ;
wire \RegFile/_1853_ ;
wire \RegFile/_1854_ ;
wire \RegFile/_1855_ ;
wire \RegFile/_1856_ ;
wire \RegFile/_1857_ ;
wire \RegFile/_1858_ ;
wire \RegFile/_1859_ ;
wire \RegFile/_1860_ ;
wire \RegFile/_1861_ ;
wire \RegFile/_1862_ ;
wire \RegFile/_1863_ ;
wire \RegFile/_1864_ ;
wire \RegFile/_1865_ ;
wire \RegFile/_1866_ ;
wire \RegFile/_1867_ ;
wire \RegFile/_1868_ ;
wire \RegFile/_1869_ ;
wire \RegFile/_1870_ ;
wire \RegFile/_1871_ ;
wire \RegFile/_1872_ ;
wire \RegFile/_1873_ ;
wire \RegFile/_1874_ ;
wire \RegFile/_1875_ ;
wire \RegFile/_1876_ ;
wire \RegFile/_1877_ ;
wire \RegFile/_1878_ ;
wire \RegFile/_1879_ ;
wire \RegFile/_1880_ ;
wire \RegFile/_1881_ ;
wire \RegFile/_1882_ ;
wire \RegFile/_1883_ ;
wire \RegFile/_1884_ ;
wire \RegFile/_1885_ ;
wire \RegFile/_1886_ ;
wire \RegFile/_1887_ ;
wire \RegFile/_1888_ ;
wire \RegFile/_1889_ ;
wire \RegFile/_1890_ ;
wire \RegFile/_1891_ ;
wire \RegFile/_1892_ ;
wire \RegFile/_1893_ ;
wire \RegFile/_1894_ ;
wire \RegFile/_1895_ ;
wire \RegFile/_1896_ ;
wire \RegFile/_1897_ ;
wire \RegFile/_1898_ ;
wire \RegFile/_1899_ ;
wire \RegFile/_1900_ ;
wire \RegFile/_1901_ ;
wire \RegFile/_1902_ ;
wire \RegFile/_1903_ ;
wire \RegFile/_1904_ ;
wire \RegFile/_1905_ ;
wire \RegFile/_1906_ ;
wire \RegFile/_1907_ ;
wire \RegFile/_1908_ ;
wire \RegFile/_1909_ ;
wire \RegFile/_1910_ ;
wire \RegFile/_1911_ ;
wire \RegFile/_1912_ ;
wire \RegFile/_1913_ ;
wire \RegFile/_1914_ ;
wire \RegFile/_1915_ ;
wire \RegFile/_1916_ ;
wire \RegFile/_1917_ ;
wire \RegFile/_1918_ ;
wire \RegFile/_1919_ ;
wire \RegFile/_1920_ ;
wire \RegFile/_1921_ ;
wire \RegFile/_1922_ ;
wire \RegFile/_1923_ ;
wire \RegFile/_1924_ ;
wire \RegFile/_1925_ ;
wire \RegFile/_1926_ ;
wire \RegFile/_1927_ ;
wire \RegFile/_1928_ ;
wire \RegFile/_1929_ ;
wire \RegFile/_1930_ ;
wire \RegFile/_1931_ ;
wire \RegFile/_1932_ ;
wire \RegFile/_1933_ ;
wire \RegFile/_1934_ ;
wire \RegFile/_1935_ ;
wire \RegFile/_1936_ ;
wire \RegFile/_1937_ ;
wire \RegFile/_1938_ ;
wire \RegFile/_1939_ ;
wire \RegFile/_1940_ ;
wire \RegFile/_1941_ ;
wire \RegFile/_1942_ ;
wire \RegFile/_1943_ ;
wire \RegFile/_1944_ ;
wire \RegFile/_1945_ ;
wire \RegFile/_1946_ ;
wire \RegFile/_1947_ ;
wire \RegFile/_1948_ ;
wire \RegFile/_1949_ ;
wire \RegFile/_1950_ ;
wire \RegFile/_1951_ ;
wire \RegFile/_1952_ ;
wire \RegFile/_1953_ ;
wire \RegFile/_1954_ ;
wire \RegFile/_1955_ ;
wire \RegFile/_1956_ ;
wire \RegFile/_1957_ ;
wire \RegFile/_1958_ ;
wire \RegFile/_1959_ ;
wire \RegFile/_1960_ ;
wire \RegFile/_1961_ ;
wire \RegFile/_1962_ ;
wire \RegFile/_1963_ ;
wire \RegFile/_1964_ ;
wire \RegFile/_1965_ ;
wire \RegFile/_1966_ ;
wire \RegFile/_1967_ ;
wire \RegFile/_1968_ ;
wire \RegFile/_1969_ ;
wire \RegFile/_1970_ ;
wire \RegFile/_1971_ ;
wire \RegFile/_1972_ ;
wire \RegFile/_1973_ ;
wire \RegFile/_1974_ ;
wire \RegFile/_1975_ ;
wire \RegFile/_1976_ ;
wire \RegFile/_1977_ ;
wire \RegFile/_1978_ ;
wire \RegFile/_1979_ ;
wire \RegFile/_1980_ ;
wire \RegFile/_1981_ ;
wire \RegFile/_1982_ ;
wire \RegFile/_1983_ ;
wire \RegFile/_1984_ ;
wire \RegFile/_1985_ ;
wire \RegFile/_1986_ ;
wire \RegFile/_1987_ ;
wire \RegFile/_1988_ ;
wire \RegFile/_1989_ ;
wire \RegFile/_1990_ ;
wire \RegFile/_1991_ ;
wire \RegFile/_1992_ ;
wire \RegFile/_1993_ ;
wire \RegFile/_1994_ ;
wire \RegFile/_1995_ ;
wire \RegFile/_1996_ ;
wire \RegFile/_1997_ ;
wire \RegFile/_1998_ ;
wire \RegFile/_1999_ ;
wire \RegFile/_2000_ ;
wire \RegFile/_2001_ ;
wire \RegFile/_2002_ ;
wire \RegFile/_2003_ ;
wire \RegFile/_2004_ ;
wire \RegFile/_2005_ ;
wire \RegFile/_2006_ ;
wire \RegFile/_2007_ ;
wire \RegFile/_2008_ ;
wire \RegFile/_2009_ ;
wire \RegFile/_2010_ ;
wire \RegFile/_2011_ ;
wire \RegFile/_2012_ ;
wire \RegFile/_2013_ ;
wire \RegFile/_2014_ ;
wire \RegFile/_2015_ ;
wire \RegFile/_2016_ ;
wire \RegFile/_2017_ ;
wire \RegFile/_2018_ ;
wire \RegFile/_2019_ ;
wire \RegFile/_2020_ ;
wire \RegFile/_2021_ ;
wire \RegFile/_2022_ ;
wire \RegFile/_2023_ ;
wire \RegFile/_2024_ ;
wire \RegFile/_2025_ ;
wire \RegFile/_2026_ ;
wire \RegFile/_2027_ ;
wire \RegFile/_2028_ ;
wire \RegFile/_2029_ ;
wire \RegFile/_2030_ ;
wire \RegFile/_2031_ ;
wire \RegFile/_2032_ ;
wire \RegFile/_2033_ ;
wire \RegFile/_2034_ ;
wire \RegFile/_2035_ ;
wire \RegFile/_2036_ ;
wire \RegFile/_2037_ ;
wire \RegFile/_2038_ ;
wire \RegFile/_2039_ ;
wire \RegFile/_2040_ ;
wire \RegFile/_2041_ ;
wire \RegFile/_2042_ ;
wire \RegFile/_2043_ ;
wire \RegFile/_2044_ ;
wire \RegFile/_2045_ ;
wire \RegFile/_2046_ ;
wire \RegFile/_2047_ ;
wire \RegFile/_2048_ ;
wire \RegFile/_2049_ ;
wire \RegFile/_2050_ ;
wire \RegFile/_2051_ ;
wire \RegFile/_2052_ ;
wire \RegFile/_2053_ ;
wire \RegFile/_2054_ ;
wire \RegFile/_2055_ ;
wire \RegFile/_2056_ ;
wire \RegFile/_2057_ ;
wire \RegFile/_2058_ ;
wire \RegFile/_2059_ ;
wire \RegFile/_2060_ ;
wire \RegFile/_2061_ ;
wire \RegFile/_2062_ ;
wire \RegFile/_2063_ ;
wire \RegFile/_2064_ ;
wire \RegFile/_2065_ ;
wire \RegFile/_2066_ ;
wire \RegFile/_2067_ ;
wire \RegFile/_2068_ ;
wire \RegFile/_2069_ ;
wire \RegFile/_2070_ ;
wire \RegFile/_2071_ ;
wire \RegFile/_2072_ ;
wire \RegFile/_2073_ ;
wire \RegFile/_2074_ ;
wire \RegFile/_2075_ ;
wire \RegFile/_2076_ ;
wire \RegFile/_2077_ ;
wire \RegFile/_2078_ ;
wire \RegFile/_2079_ ;
wire \RegFile/_2080_ ;
wire \RegFile/_2081_ ;
wire \RegFile/_2082_ ;
wire \RegFile/_2083_ ;
wire \RegFile/_2084_ ;
wire \RegFile/_2085_ ;
wire \RegFile/_2086_ ;
wire \RegFile/_2087_ ;
wire \RegFile/_2088_ ;
wire \RegFile/_2089_ ;
wire \RegFile/_2090_ ;
wire \RegFile/_2091_ ;
wire \RegFile/_2092_ ;
wire \RegFile/_2093_ ;
wire \RegFile/_2094_ ;
wire \RegFile/_2095_ ;
wire \RegFile/_2096_ ;
wire \RegFile/_2097_ ;
wire \RegFile/_2098_ ;
wire \RegFile/_2099_ ;
wire \RegFile/_2100_ ;
wire \RegFile/_2101_ ;
wire \RegFile/_2102_ ;
wire \RegFile/_2103_ ;
wire \RegFile/_2104_ ;
wire \RegFile/_2105_ ;
wire \RegFile/_2106_ ;
wire \RegFile/_2107_ ;
wire \RegFile/_2108_ ;
wire \RegFile/_2109_ ;
wire \RegFile/_2110_ ;
wire \RegFile/_2111_ ;
wire \RegFile/_2112_ ;
wire \RegFile/_2113_ ;
wire \RegFile/_2114_ ;
wire \RegFile/_2115_ ;
wire \RegFile/_2116_ ;
wire \RegFile/_2117_ ;
wire \RegFile/_2118_ ;
wire \RegFile/_2119_ ;
wire \RegFile/_2120_ ;
wire \RegFile/_2121_ ;
wire \RegFile/_2122_ ;
wire \RegFile/_2123_ ;
wire \RegFile/_2124_ ;
wire \RegFile/_2125_ ;
wire \RegFile/_2126_ ;
wire \RegFile/_2127_ ;
wire \RegFile/_2128_ ;
wire \RegFile/_2129_ ;
wire \RegFile/_2130_ ;
wire \RegFile/_2131_ ;
wire \RegFile/_2132_ ;
wire \RegFile/_2133_ ;
wire \RegFile/_2134_ ;
wire \RegFile/_2135_ ;
wire \RegFile/_2136_ ;
wire \RegFile/_2137_ ;
wire \RegFile/_2138_ ;
wire \RegFile/_2139_ ;
wire \RegFile/_2140_ ;
wire \RegFile/_2141_ ;
wire \RegFile/_2142_ ;
wire \RegFile/_2143_ ;
wire \RegFile/_2144_ ;
wire \RegFile/_2145_ ;
wire \RegFile/_2146_ ;
wire \RegFile/_2147_ ;
wire \RegFile/_2148_ ;
wire \RegFile/_2149_ ;
wire \RegFile/_2150_ ;
wire \RegFile/_2151_ ;
wire \RegFile/_2152_ ;
wire \RegFile/_2153_ ;
wire \RegFile/_2154_ ;
wire \RegFile/_2155_ ;
wire \RegFile/_2156_ ;
wire \RegFile/_2157_ ;
wire \RegFile/_2158_ ;
wire \RegFile/_2159_ ;
wire \RegFile/_2160_ ;
wire \RegFile/_2161_ ;
wire \RegFile/_2162_ ;
wire \RegFile/_2163_ ;
wire \RegFile/_2164_ ;
wire \RegFile/_2165_ ;
wire \RegFile/_2166_ ;
wire \RegFile/_2167_ ;
wire \RegFile/_2168_ ;
wire \RegFile/_2169_ ;
wire \RegFile/_2170_ ;
wire \RegFile/_2171_ ;
wire \RegFile/_2172_ ;
wire \RegFile/_2173_ ;
wire \RegFile/_2174_ ;
wire \RegFile/_2175_ ;
wire \RegFile/_2176_ ;
wire \RegFile/_2177_ ;
wire \RegFile/_2178_ ;
wire \RegFile/_2179_ ;
wire \RegFile/_2180_ ;
wire \RegFile/_2181_ ;
wire \RegFile/_2182_ ;
wire \RegFile/_2183_ ;
wire \RegFile/_2184_ ;
wire \RegFile/_2185_ ;
wire \RegFile/_2186_ ;
wire \RegFile/_2187_ ;
wire \RegFile/_2188_ ;
wire \RegFile/_2189_ ;
wire \RegFile/_2190_ ;
wire \RegFile/_2191_ ;
wire \RegFile/_2192_ ;
wire \RegFile/_2193_ ;
wire \RegFile/_2194_ ;
wire \RegFile/_2195_ ;
wire \RegFile/_2196_ ;
wire \RegFile/_2197_ ;
wire \RegFile/_2198_ ;
wire \RegFile/_2199_ ;
wire \RegFile/_2200_ ;
wire \RegFile/_2201_ ;
wire \RegFile/_2202_ ;
wire \RegFile/_2203_ ;
wire \RegFile/_2204_ ;
wire \RegFile/_2205_ ;
wire \RegFile/_2206_ ;
wire \RegFile/_2207_ ;
wire \RegFile/_2208_ ;
wire \RegFile/_2209_ ;
wire \RegFile/_2210_ ;
wire \RegFile/_2211_ ;
wire \RegFile/_2212_ ;
wire \RegFile/_2213_ ;
wire \RegFile/_2214_ ;
wire \RegFile/_2215_ ;
wire \RegFile/_2216_ ;
wire \RegFile/_2217_ ;
wire \RegFile/_2218_ ;
wire \RegFile/_2219_ ;
wire \RegFile/_2220_ ;
wire \RegFile/_2221_ ;
wire \RegFile/_2222_ ;
wire \RegFile/_2223_ ;
wire \RegFile/_2224_ ;
wire \RegFile/_2225_ ;
wire \RegFile/_2226_ ;
wire \RegFile/_2227_ ;
wire \RegFile/_2228_ ;
wire \RegFile/_2229_ ;
wire \RegFile/_2230_ ;
wire \RegFile/_2231_ ;
wire \RegFile/_2232_ ;
wire \RegFile/_2233_ ;
wire \RegFile/_2234_ ;
wire \RegFile/_2235_ ;
wire \RegFile/_2236_ ;
wire \RegFile/_2237_ ;
wire \RegFile/_2238_ ;
wire \RegFile/_2239_ ;
wire \RegFile/_2240_ ;
wire \RegFile/_2241_ ;
wire \RegFile/_2242_ ;
wire \RegFile/_2243_ ;
wire \RegFile/_2244_ ;
wire \RegFile/_2245_ ;
wire \RegFile/_2246_ ;
wire \RegFile/_2247_ ;
wire \RegFile/_2248_ ;
wire \RegFile/_2249_ ;
wire \RegFile/_2250_ ;
wire \RegFile/_2251_ ;
wire \RegFile/_2252_ ;
wire \RegFile/_2253_ ;
wire \RegFile/_2254_ ;
wire \RegFile/_2255_ ;
wire \RegFile/_2256_ ;
wire \RegFile/_2257_ ;
wire \RegFile/_2258_ ;
wire \RegFile/_2259_ ;
wire \RegFile/_2260_ ;
wire \RegFile/_2261_ ;
wire \RegFile/_2262_ ;
wire \RegFile/_2263_ ;
wire \RegFile/_2264_ ;
wire \RegFile/_2265_ ;
wire \RegFile/_2266_ ;
wire \RegFile/_2267_ ;
wire \RegFile/_2268_ ;
wire \RegFile/_2269_ ;
wire \RegFile/_2270_ ;
wire \RegFile/_2271_ ;
wire \RegFile/_2272_ ;
wire \RegFile/_2273_ ;
wire \RegFile/_2274_ ;
wire \RegFile/_2275_ ;
wire \RegFile/_2276_ ;
wire \RegFile/_2277_ ;
wire \RegFile/_2278_ ;
wire \RegFile/_2279_ ;
wire \RegFile/_2280_ ;
wire \RegFile/_2281_ ;
wire \RegFile/_2282_ ;
wire \RegFile/_2283_ ;
wire \RegFile/_2284_ ;
wire \RegFile/_2285_ ;
wire \RegFile/_2286_ ;
wire \RegFile/_2287_ ;
wire \RegFile/_2288_ ;
wire \RegFile/_2289_ ;
wire \RegFile/_2290_ ;
wire \RegFile/_2291_ ;
wire \RegFile/_2292_ ;
wire \RegFile/_2293_ ;
wire \RegFile/_2294_ ;
wire \RegFile/_2295_ ;
wire \RegFile/_2296_ ;
wire \RegFile/_2297_ ;
wire \RegFile/_2298_ ;
wire \RegFile/_2299_ ;
wire \RegFile/_2300_ ;
wire \RegFile/_2301_ ;
wire \RegFile/_2302_ ;
wire \RegFile/_2303_ ;
wire \RegFile/_2304_ ;
wire \RegFile/_2305_ ;
wire \RegFile/_2306_ ;
wire \RegFile/_2307_ ;
wire \RegFile/_2308_ ;
wire \RegFile/_2309_ ;
wire \RegFile/_2310_ ;
wire \RegFile/_2311_ ;
wire \RegFile/_2312_ ;
wire \RegFile/_2313_ ;
wire \RegFile/_2314_ ;
wire \RegFile/_2315_ ;
wire \RegFile/_2316_ ;
wire \RegFile/_2317_ ;
wire \RegFile/_2318_ ;
wire \RegFile/_2319_ ;
wire \RegFile/_2320_ ;
wire \RegFile/_2321_ ;
wire \RegFile/_2322_ ;
wire \RegFile/_2323_ ;
wire \RegFile/_2324_ ;
wire \RegFile/_2325_ ;
wire \RegFile/_2326_ ;
wire \RegFile/_2327_ ;
wire \RegFile/_2328_ ;
wire \RegFile/_2329_ ;
wire \RegFile/_2330_ ;
wire \RegFile/_2331_ ;
wire \RegFile/_2332_ ;
wire \RegFile/_2333_ ;
wire \RegFile/_2334_ ;
wire \RegFile/_2335_ ;
wire \RegFile/_2336_ ;
wire \RegFile/_2337_ ;
wire \RegFile/_2338_ ;
wire \RegFile/_2339_ ;
wire \RegFile/_2340_ ;
wire \RegFile/_2341_ ;
wire \RegFile/_2342_ ;
wire \RegFile/_2343_ ;
wire \RegFile/_2344_ ;
wire \RegFile/_2345_ ;
wire \RegFile/_2346_ ;
wire \RegFile/_2347_ ;
wire \RegFile/_2348_ ;
wire \RegFile/_2349_ ;
wire \RegFile/_2350_ ;
wire \RegFile/_2351_ ;
wire \RegFile/_2352_ ;
wire \RegFile/_2353_ ;
wire \RegFile/_2354_ ;
wire \RegFile/_2355_ ;
wire \RegFile/_2356_ ;
wire \RegFile/_2357_ ;
wire \RegFile/_2358_ ;
wire \RegFile/_2359_ ;
wire \RegFile/_2360_ ;
wire \RegFile/_2361_ ;
wire \RegFile/_2362_ ;
wire \RegFile/_2363_ ;
wire \RegFile/_2364_ ;
wire \RegFile/_2365_ ;
wire \RegFile/_2366_ ;
wire \RegFile/_2367_ ;
wire \RegFile/_2368_ ;
wire \RegFile/_2369_ ;
wire \RegFile/_2370_ ;
wire \RegFile/_2371_ ;
wire \RegFile/_2372_ ;
wire \RegFile/_2373_ ;
wire \RegFile/_2374_ ;
wire \RegFile/_2375_ ;
wire \RegFile/_2376_ ;
wire \RegFile/_2377_ ;
wire \RegFile/_2378_ ;
wire \RegFile/_2379_ ;
wire \RegFile/_2380_ ;
wire \RegFile/_2381_ ;
wire \RegFile/_2382_ ;
wire \RegFile/_2383_ ;
wire \RegFile/_2384_ ;
wire \RegFile/_2385_ ;
wire \RegFile/_2386_ ;
wire \RegFile/_2387_ ;
wire \RegFile/_2388_ ;
wire \RegFile/_2389_ ;
wire \RegFile/_2390_ ;
wire \RegFile/_2391_ ;
wire \RegFile/_2392_ ;
wire \RegFile/_2393_ ;
wire \RegFile/_2394_ ;
wire \RegFile/_2395_ ;
wire \RegFile/_2396_ ;
wire \RegFile/_2397_ ;
wire \RegFile/_2398_ ;
wire \RegFile/_2399_ ;
wire \RegFile/_2400_ ;
wire \RegFile/_2401_ ;
wire \RegFile/_2402_ ;
wire \RegFile/_2403_ ;
wire \RegFile/_2404_ ;
wire \RegFile/_2405_ ;
wire \RegFile/_2406_ ;
wire \RegFile/_2407_ ;
wire \RegFile/_2408_ ;
wire \RegFile/_2409_ ;
wire \RegFile/_2410_ ;
wire \RegFile/_2411_ ;
wire \RegFile/_2412_ ;
wire \RegFile/_2413_ ;
wire \RegFile/_2414_ ;
wire \RegFile/_2415_ ;
wire \RegFile/_2416_ ;
wire \RegFile/_2417_ ;
wire \RegFile/_2418_ ;
wire \RegFile/_2419_ ;
wire \RegFile/_2420_ ;
wire \RegFile/_2421_ ;
wire \RegFile/_2422_ ;
wire \RegFile/_2423_ ;
wire \RegFile/_2424_ ;
wire \RegFile/_2425_ ;
wire \RegFile/_2426_ ;
wire \RegFile/_2427_ ;
wire \RegFile/_2428_ ;
wire \RegFile/_2429_ ;
wire \RegFile/_2430_ ;
wire \RegFile/_2431_ ;
wire \RegFile/_2432_ ;
wire \RegFile/_2433_ ;
wire \RegFile/_2434_ ;
wire \RegFile/_2435_ ;
wire \RegFile/_2436_ ;
wire \RegFile/_2437_ ;
wire \RegFile/_2438_ ;
wire \RegFile/_2439_ ;
wire \RegFile/_2440_ ;
wire \RegFile/_2441_ ;
wire \RegFile/_2442_ ;
wire \RegFile/_2443_ ;
wire \RegFile/_2444_ ;
wire \RegFile/_2445_ ;
wire \RegFile/_2446_ ;
wire \RegFile/_2447_ ;
wire \RegFile/_2448_ ;
wire \RegFile/_2449_ ;
wire \RegFile/_2450_ ;
wire \RegFile/_2451_ ;
wire \RegFile/_2452_ ;
wire \RegFile/_2453_ ;
wire \RegFile/_2454_ ;
wire \RegFile/_2455_ ;
wire \RegFile/_2456_ ;
wire \RegFile/_2457_ ;
wire \RegFile/_2458_ ;
wire \RegFile/_2459_ ;
wire \RegFile/_2460_ ;
wire \RegFile/_2461_ ;
wire \RegFile/_2462_ ;
wire \RegFile/_2463_ ;
wire \RegFile/_2464_ ;
wire \RegFile/_2465_ ;
wire \RegFile/_2466_ ;
wire \RegFile/_2467_ ;
wire \RegFile/_2468_ ;
wire \RegFile/_2469_ ;
wire \RegFile/_2470_ ;
wire \RegFile/_2471_ ;
wire \RegFile/_2472_ ;
wire \RegFile/_2473_ ;
wire \RegFile/_2474_ ;
wire \RegFile/_2475_ ;
wire \RegFile/_2476_ ;
wire \RegFile/_2477_ ;
wire \RegFile/_2478_ ;
wire \RegFile/_2479_ ;
wire \RegFile/_2480_ ;
wire \RegFile/_2481_ ;
wire \RegFile/_2482_ ;
wire \RegFile/_2483_ ;
wire \RegFile/_2484_ ;
wire \RegFile/_2485_ ;
wire \RegFile/_2486_ ;
wire \RegFile/_2487_ ;
wire \RegFile/_2488_ ;
wire \RegFile/_2489_ ;
wire \RegFile/_2490_ ;
wire \RegFile/_2491_ ;
wire \RegFile/_2492_ ;
wire \RegFile/_2493_ ;
wire \RegFile/_2494_ ;
wire \RegFile/_2495_ ;
wire \RegFile/_2496_ ;
wire \RegFile/_2497_ ;
wire \RegFile/_2498_ ;
wire \RegFile/_2499_ ;
wire \RegFile/_2500_ ;
wire \RegFile/_2501_ ;
wire \RegFile/_2502_ ;
wire \RegFile/_2503_ ;
wire \RegFile/_2504_ ;
wire \RegFile/_2505_ ;
wire \RegFile/_2506_ ;
wire \RegFile/_2507_ ;
wire \RegFile/_2508_ ;
wire \RegFile/_2509_ ;
wire \RegFile/_2510_ ;
wire \RegFile/_2511_ ;
wire \RegFile/_2512_ ;
wire \RegFile/_2513_ ;
wire \RegFile/_2514_ ;
wire \RegFile/_2515_ ;
wire \RegFile/_2516_ ;
wire \RegFile/_2517_ ;
wire \RegFile/_2518_ ;
wire \RegFile/_2519_ ;
wire \RegFile/_2520_ ;
wire \RegFile/_2521_ ;
wire \RegFile/_2522_ ;
wire \RegFile/_2523_ ;
wire \RegFile/_2524_ ;
wire \RegFile/_2525_ ;
wire \RegFile/_2526_ ;
wire \RegFile/_2527_ ;
wire \RegFile/_2528_ ;
wire \RegFile/_2529_ ;
wire \RegFile/_2530_ ;
wire \RegFile/_2531_ ;
wire \RegFile/_2532_ ;
wire \RegFile/_2533_ ;
wire \RegFile/_2534_ ;
wire \RegFile/_2535_ ;
wire \RegFile/_2536_ ;
wire \RegFile/_2537_ ;
wire \RegFile/_2538_ ;
wire \RegFile/_2539_ ;
wire \RegFile/_2540_ ;
wire \RegFile/_2541_ ;
wire \RegFile/_2542_ ;
wire \RegFile/_2543_ ;
wire \RegFile/_2544_ ;
wire \RegFile/_2545_ ;
wire \RegFile/_2546_ ;
wire \RegFile/_2547_ ;
wire \RegFile/_2548_ ;
wire \RegFile/_2549_ ;
wire \RegFile/_2550_ ;
wire \RegFile/_2551_ ;
wire \RegFile/_2552_ ;
wire \RegFile/_2553_ ;
wire \RegFile/_2554_ ;
wire \RegFile/_2555_ ;
wire \RegFile/_2556_ ;
wire \RegFile/_2557_ ;
wire \RegFile/_2558_ ;
wire \RegFile/_2559_ ;
wire \RegFile/_2560_ ;
wire \RegFile/_2561_ ;
wire \RegFile/_2562_ ;
wire \RegFile/_2563_ ;
wire \RegFile/_2564_ ;
wire \RegFile/_2565_ ;
wire \RegFile/_2566_ ;
wire \RegFile/_2567_ ;
wire \RegFile/_2568_ ;
wire \RegFile/_2569_ ;
wire \RegFile/_2570_ ;
wire \RegFile/_2571_ ;
wire \RegFile/_2572_ ;
wire \RegFile/_2573_ ;
wire \RegFile/_2574_ ;
wire \RegFile/_2575_ ;
wire \RegFile/_2576_ ;
wire \RegFile/_2577_ ;
wire \RegFile/_2578_ ;
wire \RegFile/_2579_ ;
wire \RegFile/_2580_ ;
wire \RegFile/_2581_ ;
wire \RegFile/_2582_ ;
wire \RegFile/_2583_ ;
wire \RegFile/_2584_ ;
wire \RegFile/_2585_ ;
wire \RegFile/_2586_ ;
wire \RegFile/_2587_ ;
wire \RegFile/_2588_ ;
wire \RegFile/_2589_ ;
wire \RegFile/_2590_ ;
wire \RegFile/_2591_ ;
wire \RegFile/_2592_ ;
wire \RegFile/_2593_ ;
wire \RegFile/_2594_ ;
wire \RegFile/_2595_ ;
wire \RegFile/_2596_ ;
wire \RegFile/_2597_ ;
wire \RegFile/_2598_ ;
wire \RegFile/_2599_ ;
wire \RegFile/_2600_ ;
wire \RegFile/_2601_ ;
wire \RegFile/_2602_ ;
wire \RegFile/_2603_ ;
wire \RegFile/_2604_ ;
wire \RegFile/_2605_ ;
wire \RegFile/_2606_ ;
wire \RegFile/_2607_ ;
wire \RegFile/_2608_ ;
wire \RegFile/_2609_ ;
wire \RegFile/_2610_ ;
wire \RegFile/_2611_ ;
wire \RegFile/_2612_ ;
wire \RegFile/_2613_ ;
wire \RegFile/_2614_ ;
wire \RegFile/_2615_ ;
wire \RegFile/_2616_ ;
wire \RegFile/_2617_ ;
wire \RegFile/_2618_ ;
wire \RegFile/_2619_ ;
wire \RegFile/_2620_ ;
wire \RegFile/_2621_ ;
wire \RegFile/_2622_ ;
wire \RegFile/_2623_ ;
wire \RegFile/_2624_ ;
wire \RegFile/_2625_ ;
wire \RegFile/_2626_ ;
wire \RegFile/_2627_ ;
wire \RegFile/_2628_ ;
wire \RegFile/_2629_ ;
wire \RegFile/_2630_ ;
wire \RegFile/_2631_ ;
wire \RegFile/_2632_ ;
wire \RegFile/_2633_ ;
wire \RegFile/_2634_ ;
wire \RegFile/_2635_ ;
wire \RegFile/_2636_ ;
wire \RegFile/_2637_ ;
wire \RegFile/_2638_ ;
wire \RegFile/_2639_ ;
wire \RegFile/_2640_ ;
wire \RegFile/_2641_ ;
wire \RegFile/_2642_ ;
wire \RegFile/_2643_ ;
wire \RegFile/_2644_ ;
wire \RegFile/_2645_ ;
wire \RegFile/_2646_ ;
wire \RegFile/_2647_ ;
wire \RegFile/_2648_ ;
wire \RegFile/_2649_ ;
wire \RegFile/_2650_ ;
wire \RegFile/_2651_ ;
wire \RegFile/_2652_ ;
wire \RegFile/_2653_ ;
wire \RegFile/_2654_ ;
wire \RegFile/_2655_ ;
wire \RegFile/_2656_ ;
wire \RegFile/_2657_ ;
wire \RegFile/_2658_ ;
wire \RegFile/_2659_ ;
wire \RegFile/_2660_ ;
wire \RegFile/_2661_ ;
wire \RegFile/_2662_ ;
wire \RegFile/_2663_ ;
wire \RegFile/_2664_ ;
wire \RegFile/_2665_ ;
wire \RegFile/_2666_ ;
wire \RegFile/_2667_ ;
wire \RegFile/_2668_ ;
wire \RegFile/_2669_ ;
wire \RegFile/_2670_ ;
wire \RegFile/_2671_ ;
wire \RegFile/_2672_ ;
wire \RegFile/_2673_ ;
wire \RegFile/_2674_ ;
wire \RegFile/_2675_ ;
wire \RegFile/_2676_ ;
wire \RegFile/_2677_ ;
wire \RegFile/_2678_ ;
wire \RegFile/_2679_ ;
wire \RegFile/_2680_ ;
wire \RegFile/_2681_ ;
wire \RegFile/_2682_ ;
wire \RegFile/_2683_ ;
wire \RegFile/_2684_ ;
wire \RegFile/_2685_ ;
wire \RegFile/_2686_ ;
wire \RegFile/_2687_ ;
wire \RegFile/_2688_ ;
wire \RegFile/_2689_ ;
wire \RegFile/_2690_ ;
wire \RegFile/_2691_ ;
wire \RegFile/_2692_ ;
wire \RegFile/_2693_ ;
wire \RegFile/_2694_ ;
wire \RegFile/_2695_ ;
wire \RegFile/_2696_ ;
wire \RegFile/_2697_ ;
wire \RegFile/_2698_ ;
wire \RegFile/_2699_ ;
wire \RegFile/_2700_ ;
wire \RegFile/_2701_ ;
wire \RegFile/_2702_ ;
wire \RegFile/_2703_ ;
wire \RegFile/_2704_ ;
wire \RegFile/_2705_ ;
wire \RegFile/_2706_ ;
wire \RegFile/_2707_ ;
wire \RegFile/_2708_ ;
wire \RegFile/_2709_ ;
wire \RegFile/_2710_ ;
wire \RegFile/_2711_ ;
wire \RegFile/_2712_ ;
wire \RegFile/_2713_ ;
wire \RegFile/_2714_ ;
wire \RegFile/_2715_ ;
wire \RegFile/_2716_ ;
wire \RegFile/_2717_ ;
wire \RegFile/_2718_ ;
wire \RegFile/_2719_ ;
wire \RegFile/_2720_ ;
wire \RegFile/_2721_ ;
wire \RegFile/_2722_ ;
wire \RegFile/_2723_ ;
wire \RegFile/_2724_ ;
wire \RegFile/_2725_ ;
wire \RegFile/_2726_ ;
wire \RegFile/_2727_ ;
wire \RegFile/_2728_ ;
wire \RegFile/_2729_ ;
wire \RegFile/_2730_ ;
wire \RegFile/_2731_ ;
wire \RegFile/_2732_ ;
wire \RegFile/_2733_ ;
wire \RegFile/_2734_ ;
wire \RegFile/_2735_ ;
wire \RegFile/_2736_ ;
wire \RegFile/_2737_ ;
wire \RegFile/_2738_ ;
wire \RegFile/_2739_ ;
wire \RegFile/_2740_ ;
wire \RegFile/_2741_ ;
wire \RegFile/_2742_ ;
wire \RegFile/_2743_ ;
wire \RegFile/_2744_ ;
wire \RegFile/_2745_ ;
wire \RegFile/_2746_ ;
wire \RegFile/_2747_ ;
wire \RegFile/_2748_ ;
wire \RegFile/_2749_ ;
wire \RegFile/_2750_ ;
wire \RegFile/_2751_ ;
wire \RegFile/_2752_ ;
wire \RegFile/_2753_ ;
wire \RegFile/_2754_ ;
wire \RegFile/_2755_ ;
wire \RegFile/_2756_ ;
wire \RegFile/_2757_ ;
wire \RegFile/_2758_ ;
wire \RegFile/_2759_ ;
wire \RegFile/_2760_ ;
wire \RegFile/_2761_ ;
wire \RegFile/_2762_ ;
wire \RegFile/_2763_ ;
wire \RegFile/_2764_ ;
wire \RegFile/_2765_ ;
wire \RegFile/_2766_ ;
wire \RegFile/_2767_ ;
wire \RegFile/_2768_ ;
wire \RegFile/_2769_ ;
wire \RegFile/_2770_ ;
wire \RegFile/_2771_ ;
wire \RegFile/_2772_ ;
wire \RegFile/_2773_ ;
wire \RegFile/_2774_ ;
wire \RegFile/_2775_ ;
wire \RegFile/_2776_ ;
wire \RegFile/_2777_ ;
wire \RegFile/_2778_ ;
wire \RegFile/_2779_ ;
wire \RegFile/_2780_ ;
wire \RegFile/_2781_ ;
wire \RegFile/_2782_ ;
wire \RegFile/_2783_ ;
wire \RegFile/_2784_ ;
wire \RegFile/_2785_ ;
wire \RegFile/_2786_ ;
wire \RegFile/_2787_ ;
wire \RegFile/_2788_ ;
wire \RegFile/_2789_ ;
wire \RegFile/_2790_ ;
wire \RegFile/_2791_ ;
wire \RegFile/_2792_ ;
wire \RegFile/_2793_ ;
wire \RegFile/_2794_ ;
wire \RegFile/_2795_ ;
wire \RegFile/_2796_ ;
wire \RegFile/_2797_ ;
wire \RegFile/_2798_ ;
wire \RegFile/_2799_ ;
wire \RegFile/_2800_ ;
wire \RegFile/_2801_ ;
wire \RegFile/_2802_ ;
wire \RegFile/_2803_ ;
wire \RegFile/_2804_ ;
wire \RegFile/_2805_ ;
wire \RegFile/_2806_ ;
wire \RegFile/_2807_ ;
wire \RegFile/_2808_ ;
wire \RegFile/_2809_ ;
wire \RegFile/_2810_ ;
wire \RegFile/_2811_ ;
wire \RegFile/_2812_ ;
wire \RegFile/_2813_ ;
wire \RegFile/_2814_ ;
wire \RegFile/_2815_ ;
wire \RegFile/_2816_ ;
wire \RegFile/_2817_ ;
wire \RegFile/_2818_ ;
wire \RegFile/_2819_ ;
wire \RegFile/_2820_ ;
wire \RegFile/_2821_ ;
wire \RegFile/_2822_ ;
wire \RegFile/_2823_ ;
wire \RegFile/_2824_ ;
wire \RegFile/_2825_ ;
wire \RegFile/_2826_ ;
wire \RegFile/_2827_ ;
wire \RegFile/_2828_ ;
wire \RegFile/_2829_ ;
wire \RegFile/_2830_ ;
wire \RegFile/_2831_ ;
wire \RegFile/_2832_ ;
wire \RegFile/_2833_ ;
wire \RegFile/_2834_ ;
wire \RegFile/_2835_ ;
wire \RegFile/_2836_ ;
wire \RegFile/_2837_ ;
wire \RegFile/_2838_ ;
wire \RegFile/_2839_ ;
wire \RegFile/_2840_ ;
wire \RegFile/_2841_ ;
wire \RegFile/_2842_ ;
wire \RegFile/_2843_ ;
wire \RegFile/_2844_ ;
wire \RegFile/_2845_ ;
wire \RegFile/_2846_ ;
wire \RegFile/_2847_ ;
wire \RegFile/_2848_ ;
wire \RegFile/_2849_ ;
wire \RegFile/_2850_ ;
wire \RegFile/_2851_ ;
wire \RegFile/_2852_ ;
wire \RegFile/_2853_ ;
wire \RegFile/_2854_ ;
wire \RegFile/_2855_ ;
wire \RegFile/_2856_ ;
wire \RegFile/_2857_ ;
wire \RegFile/_2858_ ;
wire \RegFile/_2859_ ;
wire \RegFile/_2860_ ;
wire \RegFile/_2861_ ;
wire \RegFile/_2862_ ;
wire \RegFile/_2863_ ;
wire \RegFile/_2864_ ;
wire \RegFile/_2865_ ;
wire \RegFile/_2866_ ;
wire \RegFile/_2867_ ;
wire \RegFile/_2868_ ;
wire \RegFile/_2869_ ;
wire \RegFile/_2870_ ;
wire \RegFile/_2871_ ;
wire \RegFile/_2872_ ;
wire \RegFile/_2873_ ;
wire \RegFile/_2874_ ;
wire \RegFile/_2875_ ;
wire \RegFile/_2876_ ;
wire \RegFile/_2877_ ;
wire \RegFile/_2878_ ;
wire \RegFile/_2879_ ;
wire \RegFile/_2880_ ;
wire \RegFile/_2881_ ;
wire \RegFile/_2882_ ;
wire \RegFile/_2883_ ;
wire \RegFile/_2884_ ;
wire \RegFile/_2885_ ;
wire \RegFile/_2886_ ;
wire \RegFile/_2887_ ;
wire \RegFile/_2888_ ;
wire \RegFile/_2889_ ;
wire \RegFile/_2890_ ;
wire \RegFile/_2891_ ;
wire \RegFile/_2892_ ;
wire \RegFile/_2893_ ;
wire \RegFile/_2894_ ;
wire \RegFile/_2895_ ;
wire \RegFile/_2896_ ;
wire \RegFile/_2897_ ;
wire \RegFile/_2898_ ;
wire \RegFile/_2899_ ;
wire \RegFile/_2900_ ;
wire \RegFile/_2901_ ;
wire \RegFile/_2902_ ;
wire \RegFile/_2903_ ;
wire \RegFile/_2904_ ;
wire \RegFile/_2905_ ;
wire \RegFile/_2906_ ;
wire \RegFile/_2907_ ;
wire \RegFile/_2908_ ;
wire \RegFile/_2909_ ;
wire \RegFile/_2910_ ;
wire \RegFile/_2911_ ;
wire \RegFile/_2912_ ;
wire \RegFile/_2913_ ;
wire \RegFile/_2914_ ;
wire \RegFile/_2915_ ;
wire \RegFile/_2916_ ;
wire \RegFile/_2917_ ;
wire \RegFile/_2918_ ;
wire \RegFile/_2919_ ;
wire \RegFile/_2920_ ;
wire \RegFile/_2921_ ;
wire \RegFile/_2922_ ;
wire \RegFile/_2923_ ;
wire \RegFile/_2924_ ;
wire \RegFile/_2925_ ;
wire \RegFile/_2926_ ;
wire \RegFile/_2927_ ;
wire \RegFile/_2928_ ;
wire \RegFile/_2929_ ;
wire \RegFile/_2930_ ;
wire \RegFile/_2931_ ;
wire \RegFile/_2932_ ;
wire \RegFile/_2933_ ;
wire \RegFile/_2934_ ;
wire \RegFile/_2935_ ;
wire \RegFile/_2936_ ;
wire \RegFile/_2937_ ;
wire \RegFile/_2938_ ;
wire \RegFile/_2939_ ;
wire \RegFile/_2940_ ;
wire \RegFile/_2941_ ;
wire \RegFile/_2942_ ;
wire \RegFile/_2943_ ;
wire \RegFile/_2944_ ;
wire \RegFile/_2945_ ;
wire \RegFile/_2946_ ;
wire \RegFile/_2947_ ;
wire \RegFile/_2948_ ;
wire \RegFile/_2949_ ;
wire \RegFile/_2950_ ;
wire \RegFile/_2951_ ;
wire \RegFile/_2952_ ;
wire \RegFile/_2953_ ;
wire \RegFile/_2954_ ;
wire \RegFile/_2955_ ;
wire \RegFile/_2956_ ;
wire \RegFile/_2957_ ;
wire \RegFile/_2958_ ;
wire \RegFile/_2959_ ;
wire \RegFile/_2960_ ;
wire \RegFile/_2961_ ;
wire \RegFile/_2962_ ;
wire \RegFile/_2963_ ;
wire \RegFile/_2964_ ;
wire \RegFile/_2965_ ;
wire \RegFile/_2966_ ;
wire \RegFile/_2967_ ;
wire \RegFile/_2968_ ;
wire \RegFile/_2969_ ;
wire \RegFile/_2970_ ;
wire \RegFile/_2971_ ;
wire \RegFile/_2972_ ;
wire \RegFile/_2973_ ;
wire \RegFile/_2974_ ;
wire \RegFile/_2975_ ;
wire \RegFile/_2976_ ;
wire \RegFile/_2977_ ;
wire \RegFile/_2978_ ;
wire \RegFile/_2979_ ;
wire \RegFile/_2980_ ;
wire \RegFile/_2981_ ;
wire \RegFile/_2982_ ;
wire \RegFile/_2983_ ;
wire \RegFile/_2984_ ;
wire \RegFile/_2985_ ;
wire \RegFile/_2986_ ;
wire \RegFile/_2987_ ;
wire \RegFile/_2988_ ;
wire \RegFile/_2989_ ;
wire \RegFile/_2990_ ;
wire \RegFile/_2991_ ;
wire \RegFile/_2992_ ;
wire \RegFile/_2993_ ;
wire \RegFile/_2994_ ;
wire \RegFile/_2995_ ;
wire \RegFile/_2996_ ;
wire \RegFile/_2997_ ;
wire \RegFile/_2998_ ;
wire \RegFile/_2999_ ;
wire \RegFile/_3000_ ;
wire \RegFile/_3001_ ;
wire \RegFile/_3002_ ;
wire \RegFile/_3003_ ;
wire \RegFile/_3004_ ;
wire \RegFile/_3005_ ;
wire \RegFile/_3006_ ;
wire \RegFile/_3007_ ;
wire \RegFile/_3008_ ;
wire \RegFile/_3009_ ;
wire \RegFile/_3010_ ;
wire \RegFile/_3011_ ;
wire \RegFile/_3012_ ;
wire \RegFile/_3013_ ;
wire \RegFile/_3014_ ;
wire \RegFile/_3015_ ;
wire \RegFile/_3016_ ;
wire \RegFile/_3017_ ;
wire \RegFile/_3018_ ;
wire \RegFile/_3019_ ;
wire \RegFile/_3020_ ;
wire \RegFile/_3021_ ;
wire \RegFile/_3022_ ;
wire \RegFile/_3023_ ;
wire \RegFile/_3024_ ;
wire \RegFile/_3025_ ;
wire \RegFile/_3026_ ;
wire \RegFile/_3027_ ;
wire \RegFile/_3028_ ;
wire \RegFile/_3029_ ;
wire \RegFile/_3030_ ;
wire \RegFile/_3031_ ;
wire \RegFile/_3032_ ;
wire \RegFile/_3033_ ;
wire \RegFile/_3034_ ;
wire \RegFile/_3035_ ;
wire \RegFile/_3036_ ;
wire \RegFile/_3037_ ;
wire \RegFile/_3038_ ;
wire \RegFile/_3039_ ;
wire \RegFile/_3040_ ;
wire \RegFile/_3041_ ;
wire \RegFile/_3042_ ;
wire \RegFile/_3043_ ;
wire \RegFile/_3044_ ;
wire \RegFile/_3045_ ;
wire \RegFile/_3046_ ;
wire \RegFile/_3047_ ;
wire \RegFile/_3048_ ;
wire \RegFile/_3049_ ;
wire \RegFile/_3050_ ;
wire \RegFile/_3051_ ;
wire \RegFile/_3052_ ;
wire \RegFile/_3053_ ;
wire \RegFile/_3054_ ;
wire \RegFile/_3055_ ;
wire \RegFile/_3056_ ;
wire \RegFile/_3057_ ;
wire \RegFile/_3058_ ;
wire \RegFile/_3059_ ;
wire \RegFile/_3060_ ;
wire \RegFile/_3061_ ;
wire \RegFile/_3062_ ;
wire \RegFile/_3063_ ;
wire \RegFile/_3064_ ;
wire \RegFile/_3065_ ;
wire \RegFile/_3066_ ;
wire \RegFile/_3067_ ;
wire \RegFile/_3068_ ;
wire \RegFile/_3069_ ;
wire \RegFile/_3070_ ;
wire \RegFile/_3071_ ;
wire \RegFile/_3072_ ;
wire \RegFile/_3073_ ;
wire \RegFile/_3074_ ;
wire \RegFile/_3075_ ;
wire \RegFile/_3076_ ;
wire \RegFile/_3077_ ;
wire \RegFile/_3078_ ;
wire \RegFile/_3079_ ;
wire \RegFile/_3080_ ;
wire \RegFile/_3081_ ;
wire \RegFile/_3082_ ;
wire \RegFile/_3083_ ;
wire \RegFile/_3084_ ;
wire \RegFile/_3085_ ;
wire \RegFile/_3086_ ;
wire \RegFile/_3087_ ;
wire \RegFile/_3088_ ;
wire \RegFile/_3089_ ;
wire \RegFile/_3090_ ;
wire \RegFile/_3091_ ;
wire \RegFile/_3092_ ;
wire \RegFile/_3093_ ;
wire \RegFile/_3094_ ;
wire \RegFile/_3095_ ;
wire \RegFile/_3096_ ;
wire \RegFile/_3097_ ;
wire \RegFile/_3098_ ;
wire \RegFile/_3099_ ;
wire \RegFile/_3100_ ;
wire \RegFile/_3101_ ;
wire \RegFile/_3102_ ;
wire \RegFile/_3103_ ;
wire \RegFile/_3104_ ;
wire \RegFile/_3105_ ;
wire \RegFile/_3106_ ;
wire \RegFile/_3107_ ;
wire \RegFile/_3108_ ;
wire \RegFile/_3109_ ;
wire \RegFile/_3110_ ;
wire \RegFile/_3111_ ;
wire \RegFile/_3112_ ;
wire \RegFile/_3113_ ;
wire \RegFile/_3114_ ;
wire \RegFile/_3115_ ;
wire \RegFile/_3116_ ;
wire \RegFile/_3117_ ;
wire \RegFile/_3118_ ;
wire \RegFile/_3119_ ;
wire \RegFile/_3120_ ;
wire \RegFile/_3121_ ;
wire \RegFile/_3122_ ;
wire \RegFile/_3123_ ;
wire \RegFile/_3124_ ;
wire \RegFile/_3125_ ;
wire \RegFile/_3126_ ;
wire \RegFile/_3127_ ;
wire \RegFile/_3128_ ;
wire \RegFile/_3129_ ;
wire \RegFile/_3130_ ;
wire \RegFile/_3131_ ;
wire \RegFile/_3132_ ;
wire \RegFile/_3133_ ;
wire \RegFile/_3134_ ;
wire \RegFile/_3135_ ;
wire \RegFile/_3136_ ;
wire \RegFile/_3137_ ;
wire \RegFile/_3138_ ;
wire \RegFile/_3139_ ;
wire \RegFile/_3140_ ;
wire \RegFile/_3141_ ;
wire \RegFile/_3142_ ;
wire \RegFile/_3143_ ;
wire \RegFile/_3144_ ;
wire \RegFile/_3145_ ;
wire \RegFile/_3146_ ;
wire \RegFile/_3147_ ;
wire \RegFile/_3148_ ;
wire \RegFile/_3149_ ;
wire \RegFile/_3150_ ;
wire \RegFile/_3151_ ;
wire \RegFile/_3152_ ;
wire \RegFile/_3153_ ;
wire \RegFile/_3154_ ;
wire \RegFile/_3155_ ;
wire \RegFile/_3156_ ;
wire \RegFile/_3157_ ;
wire \RegFile/_3158_ ;
wire \RegFile/_3159_ ;
wire \RegFile/_3160_ ;
wire \RegFile/_3161_ ;
wire \RegFile/_3162_ ;
wire \RegFile/_3163_ ;
wire \RegFile/_3164_ ;
wire \RegFile/_3165_ ;
wire \RegFile/_3166_ ;
wire \RegFile/_3167_ ;
wire \RegFile/_3168_ ;
wire \RegFile/_3169_ ;
wire \RegFile/_3170_ ;
wire \RegFile/_3171_ ;
wire \RegFile/_3172_ ;
wire \RegFile/_3173_ ;
wire \RegFile/_3174_ ;
wire \RegFile/_3175_ ;
wire \RegFile/_3176_ ;
wire \RegFile/_3177_ ;
wire \RegFile/_3178_ ;
wire \RegFile/_3179_ ;
wire \RegFile/_3180_ ;
wire \RegFile/_3181_ ;
wire \RegFile/_3182_ ;
wire \RegFile/_3183_ ;
wire \RegFile/_3184_ ;
wire \RegFile/_3185_ ;
wire \RegFile/_3186_ ;
wire \RegFile/_3187_ ;
wire \RegFile/_3188_ ;
wire \RegFile/_3189_ ;
wire \RegFile/_3190_ ;
wire \RegFile/_3191_ ;
wire \RegFile/_3192_ ;
wire \RegFile/_3193_ ;
wire \RegFile/_3194_ ;
wire \RegFile/_3195_ ;
wire \RegFile/_3196_ ;
wire \RegFile/_3197_ ;
wire \RegFile/_3198_ ;
wire \RegFile/_3199_ ;
wire \RegFile/_3200_ ;
wire \RegFile/_3201_ ;
wire \RegFile/_3202_ ;
wire \RegFile/_3203_ ;
wire \RegFile/_3204_ ;
wire \RegFile/_3205_ ;
wire \RegFile/_3206_ ;
wire \RegFile/_3207_ ;
wire \RegFile/_3208_ ;
wire \RegFile/_3209_ ;
wire \RegFile/_3210_ ;
wire \RegFile/_3211_ ;
wire \RegFile/_3212_ ;
wire \RegFile/_3213_ ;
wire \RegFile/_3214_ ;
wire \RegFile/_3215_ ;
wire \RegFile/_3216_ ;
wire \RegFile/_3217_ ;
wire \RegFile/_3218_ ;
wire \RegFile/_3219_ ;
wire \RegFile/_3220_ ;
wire \RegFile/_3221_ ;
wire \RegFile/_3222_ ;
wire \RegFile/_3223_ ;
wire \RegFile/_3224_ ;
wire \RegFile/_3225_ ;
wire \RegFile/_3226_ ;
wire \RegFile/_3227_ ;
wire \RegFile/_3228_ ;
wire \RegFile/_3229_ ;
wire \RegFile/_3230_ ;
wire \RegFile/_3231_ ;
wire \RegFile/_3232_ ;
wire \RegFile/_3233_ ;
wire \RegFile/_3234_ ;
wire \RegFile/_3235_ ;
wire \RegFile/_3236_ ;
wire \RegFile/_3237_ ;
wire \RegFile/_3238_ ;
wire \RegFile/_3239_ ;
wire \RegFile/_3240_ ;
wire \RegFile/_3241_ ;
wire \RegFile/_3242_ ;
wire \RegFile/_3243_ ;
wire \RegFile/_3244_ ;
wire \RegFile/_3245_ ;
wire \RegFile/_3246_ ;
wire \RegFile/_3247_ ;
wire \RegFile/_3248_ ;
wire \RegFile/_3249_ ;
wire \RegFile/_3250_ ;
wire \RegFile/_3251_ ;
wire \RegFile/_3252_ ;
wire \RegFile/_3253_ ;
wire \RegFile/_3254_ ;
wire \RegFile/_3255_ ;
wire \RegFile/_3256_ ;
wire \RegFile/_3257_ ;
wire \RegFile/_3258_ ;
wire \RegFile/_3259_ ;
wire \RegFile/_3260_ ;
wire \RegFile/_3261_ ;
wire \RegFile/_3262_ ;
wire \RegFile/_3263_ ;
wire \RegFile/_3264_ ;
wire \RegFile/_3265_ ;
wire \RegFile/_3266_ ;
wire \RegFile/_3267_ ;
wire \RegFile/_3268_ ;
wire \RegFile/_3269_ ;
wire \RegFile/_3270_ ;
wire \RegFile/_3271_ ;
wire \RegFile/_3272_ ;
wire \RegFile/_3273_ ;
wire \RegFile/_3274_ ;
wire \RegFile/_3275_ ;
wire \RegFile/_3276_ ;
wire \RegFile/_3277_ ;
wire \RegFile/_3278_ ;
wire \RegFile/_3279_ ;
wire \RegFile/_3280_ ;
wire \RegFile/_3281_ ;
wire \RegFile/_3282_ ;
wire \RegFile/_3283_ ;
wire \RegFile/_3284_ ;
wire \RegFile/_3285_ ;
wire \RegFile/_3286_ ;
wire \RegFile/_3287_ ;
wire \RegFile/_3288_ ;
wire \RegFile/_3289_ ;
wire \RegFile/_3290_ ;
wire \RegFile/_3291_ ;
wire \RegFile/_3292_ ;
wire \RegFile/_3293_ ;
wire \RegFile/_3294_ ;
wire \RegFile/_3295_ ;
wire \RegFile/_3296_ ;
wire \RegFile/_3297_ ;
wire \RegFile/_3298_ ;
wire \RegFile/_3299_ ;
wire \RegFile/_3300_ ;
wire \RegFile/_3301_ ;
wire \RegFile/_3302_ ;
wire \RegFile/_3303_ ;
wire \RegFile/_3304_ ;
wire \RegFile/_3305_ ;
wire \RegFile/_3306_ ;
wire \RegFile/_3307_ ;
wire \RegFile/_3308_ ;
wire \RegFile/_3309_ ;
wire \RegFile/_3310_ ;
wire \RegFile/_3311_ ;
wire \RegFile/_3312_ ;
wire \RegFile/_3313_ ;
wire \RegFile/_3314_ ;
wire \RegFile/_3315_ ;
wire \RegFile/_3316_ ;
wire \RegFile/_3317_ ;
wire \RegFile/_3318_ ;
wire \RegFile/_3319_ ;
wire \RegFile/_3320_ ;
wire \RegFile/_3321_ ;
wire \RegFile/_3322_ ;
wire \RegFile/_3323_ ;
wire \RegFile/_3324_ ;
wire \RegFile/_3325_ ;
wire \RegFile/_3326_ ;
wire \RegFile/_3327_ ;
wire \RegFile/_3328_ ;
wire \RegFile/_3329_ ;
wire \RegFile/_3330_ ;
wire \RegFile/_3331_ ;
wire \RegFile/_3332_ ;
wire \RegFile/_3333_ ;
wire \RegFile/_3334_ ;
wire \RegFile/_3335_ ;
wire \RegFile/_3336_ ;
wire \RegFile/_3337_ ;
wire \RegFile/_3338_ ;
wire \RegFile/_3339_ ;
wire \RegFile/_3340_ ;
wire \RegFile/_3341_ ;
wire \RegFile/_3342_ ;
wire \RegFile/_3343_ ;
wire \RegFile/_3344_ ;
wire \RegFile/_3345_ ;
wire \RegFile/_3346_ ;
wire \RegFile/_3347_ ;
wire \RegFile/_3348_ ;
wire \RegFile/_3349_ ;
wire \RegFile/_3350_ ;
wire \RegFile/_3351_ ;
wire \RegFile/_3352_ ;
wire \RegFile/_3353_ ;
wire \RegFile/_3354_ ;
wire \RegFile/_3355_ ;
wire \RegFile/_3356_ ;
wire \RegFile/_3357_ ;
wire \RegFile/_3358_ ;
wire \RegFile/_3359_ ;
wire \RegFile/_3360_ ;
wire \RegFile/_3361_ ;
wire \RegFile/_3362_ ;
wire \RegFile/_3363_ ;
wire \RegFile/_3364_ ;
wire \RegFile/_3365_ ;
wire \RegFile/_3366_ ;
wire \RegFile/_3367_ ;
wire \RegFile/_3368_ ;
wire \RegFile/_3369_ ;
wire \RegFile/_3370_ ;
wire \RegFile/_3371_ ;
wire \RegFile/_3372_ ;
wire \RegFile/_3373_ ;
wire \RegFile/_3374_ ;
wire \RegFile/_3375_ ;
wire \RegFile/_3376_ ;
wire \RegFile/_3377_ ;
wire \RegFile/_3378_ ;
wire \RegFile/_3379_ ;
wire \RegFile/_3380_ ;
wire \RegFile/_3381_ ;
wire \RegFile/_3382_ ;
wire \RegFile/_3383_ ;
wire \RegFile/_3384_ ;
wire \RegFile/_3385_ ;
wire \RegFile/_3386_ ;
wire \RegFile/_3387_ ;
wire \RegFile/_3388_ ;
wire \RegFile/_3389_ ;
wire \RegFile/_3390_ ;
wire \RegFile/_3391_ ;
wire \RegFile/_3392_ ;
wire \RegFile/_3393_ ;
wire \RegFile/_3394_ ;
wire \RegFile/_3395_ ;
wire \RegFile/_3396_ ;
wire \RegFile/_3397_ ;
wire \RegFile/_3398_ ;
wire \RegFile/_3399_ ;
wire \RegFile/_3400_ ;
wire \RegFile/_3401_ ;
wire \RegFile/_3402_ ;
wire \RegFile/_3403_ ;
wire \RegFile/_3404_ ;
wire \RegFile/_3405_ ;
wire \RegFile/_3406_ ;
wire \RegFile/_3407_ ;
wire \RegFile/_3408_ ;
wire \RegFile/_3409_ ;
wire \RegFile/_3410_ ;
wire \RegFile/_3411_ ;
wire \RegFile/_3412_ ;
wire \RegFile/_3413_ ;
wire \RegFile/_3414_ ;
wire \RegFile/_3415_ ;
wire \RegFile/_3416_ ;
wire \RegFile/_3417_ ;
wire \RegFile/_3418_ ;
wire \RegFile/_3419_ ;
wire \RegFile/_3420_ ;
wire \RegFile/_3421_ ;
wire \RegFile/_3422_ ;
wire \RegFile/_3423_ ;
wire \RegFile/_3424_ ;
wire \RegFile/_3425_ ;
wire \RegFile/_3426_ ;
wire \RegFile/_3427_ ;
wire \RegFile/_3428_ ;
wire \RegFile/_3429_ ;
wire \RegFile/_3430_ ;
wire \RegFile/_3431_ ;
wire \RegFile/_3432_ ;
wire \RegFile/_3433_ ;
wire \RegFile/_3434_ ;
wire \RegFile/_3435_ ;
wire \RegFile/_3436_ ;
wire \RegFile/_3437_ ;
wire \RegFile/_3438_ ;
wire \RegFile/_3439_ ;
wire \RegFile/_3440_ ;
wire \RegFile/_3441_ ;
wire \RegFile/_3442_ ;
wire \RegFile/_3443_ ;
wire \RegFile/_3444_ ;
wire \RegFile/_3445_ ;
wire \RegFile/_3446_ ;
wire \RegFile/_3447_ ;
wire \RegFile/_3448_ ;
wire \RegFile/_3449_ ;
wire \RegFile/_3450_ ;
wire \RegFile/_3451_ ;
wire \RegFile/_3452_ ;
wire \RegFile/_3453_ ;
wire \RegFile/_3454_ ;
wire \RegFile/_3455_ ;
wire \RegFile/_3456_ ;
wire \RegFile/_3457_ ;
wire \RegFile/_3458_ ;
wire \RegFile/_3459_ ;
wire \RegFile/_3460_ ;
wire \RegFile/_3461_ ;
wire \RegFile/_3462_ ;
wire \RegFile/_3463_ ;
wire \RegFile/_3464_ ;
wire \RegFile/_3465_ ;
wire \RegFile/_3466_ ;
wire \RegFile/_3467_ ;
wire \RegFile/_3468_ ;
wire \RegFile/_3469_ ;
wire \RegFile/_3470_ ;
wire \RegFile/_3471_ ;
wire \RegFile/_3472_ ;
wire \RegFile/_3473_ ;
wire \RegFile/_3474_ ;
wire \RegFile/_3475_ ;
wire \RegFile/_3476_ ;
wire \RegFile/_3477_ ;
wire \RegFile/_3478_ ;
wire \RegFile/_3479_ ;
wire \RegFile/_3480_ ;
wire \RegFile/_3481_ ;
wire \RegFile/_3482_ ;
wire \RegFile/_3483_ ;
wire \RegFile/_3484_ ;
wire \RegFile/_3485_ ;
wire \RegFile/_3486_ ;
wire \RegFile/_3487_ ;
wire \RegFile/_3488_ ;
wire \RegFile/_3489_ ;
wire \RegFile/_3490_ ;
wire \RegFile/_3491_ ;
wire \RegFile/_3492_ ;
wire \RegFile/_3493_ ;
wire \RegFile/_3494_ ;
wire \RegFile/_3495_ ;
wire \RegFile/_3496_ ;
wire \RegFile/_3497_ ;
wire \RegFile/_3498_ ;
wire \RegFile/_3499_ ;
wire \RegFile/_3500_ ;
wire \RegFile/_3501_ ;
wire \RegFile/_3502_ ;
wire \RegFile/_3503_ ;
wire \RegFile/_3504_ ;
wire \RegFile/_3505_ ;
wire \RegFile/_3506_ ;
wire \RegFile/_3507_ ;
wire \RegFile/_3508_ ;
wire \RegFile/_3509_ ;
wire \RegFile/_3510_ ;
wire \RegFile/_3511_ ;
wire \RegFile/_3512_ ;
wire \RegFile/_3513_ ;
wire \RegFile/_3514_ ;
wire \RegFile/_3515_ ;
wire \RegFile/_3516_ ;
wire \RegFile/_3517_ ;
wire \RegFile/_3518_ ;
wire \RegFile/_3519_ ;
wire \RegFile/_3520_ ;
wire \RegFile/_3521_ ;
wire \RegFile/_3522_ ;
wire \RegFile/_3523_ ;
wire \RegFile/_3524_ ;
wire \RegFile/_3525_ ;
wire \RegFile/_3526_ ;
wire \RegFile/_3527_ ;
wire \RegFile/_3528_ ;
wire \RegFile/_3529_ ;
wire \RegFile/_3530_ ;
wire \RegFile/_3531_ ;
wire \RegFile/_3532_ ;
wire \RegFile/_3533_ ;
wire \RegFile/_3534_ ;
wire \RegFile/_3535_ ;
wire \RegFile/_3536_ ;
wire \RegFile/_3537_ ;
wire \RegFile/_3538_ ;
wire \RegFile/_3539_ ;
wire \RegFile/_3540_ ;
wire \RegFile/_3541_ ;
wire \RegFile/_3542_ ;
wire \RegFile/_3543_ ;
wire \RegFile/_3544_ ;
wire \RegFile/_3545_ ;
wire \RegFile/_3546_ ;
wire \RegFile/_3547_ ;
wire \RegFile/_3548_ ;
wire \RegFile/_3549_ ;
wire \RegFile/_3550_ ;
wire \RegFile/_3551_ ;
wire \RegFile/_3552_ ;
wire \RegFile/_3553_ ;
wire \RegFile/_3554_ ;
wire \RegFile/_3555_ ;
wire \RegFile/_3556_ ;
wire \RegFile/_3557_ ;
wire \RegFile/_3558_ ;
wire \RegFile/_3559_ ;
wire \RegFile/_3560_ ;
wire \RegFile/_3561_ ;
wire \RegFile/_3562_ ;
wire \RegFile/_3563_ ;
wire \RegFile/_3564_ ;
wire \RegFile/_3565_ ;
wire \RegFile/_3566_ ;
wire \RegFile/_3567_ ;
wire \RegFile/_3568_ ;
wire \RegFile/_3569_ ;
wire \RegFile/_3570_ ;
wire \RegFile/_3571_ ;
wire \RegFile/_3572_ ;
wire \RegFile/_3573_ ;
wire \RegFile/_3574_ ;
wire \RegFile/_3575_ ;
wire \RegFile/_3576_ ;
wire \RegFile/_3577_ ;
wire \RegFile/_3578_ ;
wire \RegFile/_3579_ ;
wire \RegFile/_3580_ ;
wire \RegFile/_3581_ ;
wire \RegFile/_3582_ ;
wire \RegFile/_3583_ ;
wire \RegFile/_3584_ ;
wire \RegFile/_3585_ ;
wire \RegFile/_3586_ ;
wire \RegFile/_3587_ ;
wire \RegFile/_3588_ ;
wire \RegFile/_3589_ ;
wire \RegFile/_3590_ ;
wire \RegFile/_3591_ ;
wire \RegFile/_3592_ ;
wire \RegFile/_3593_ ;
wire \RegFile/_3594_ ;
wire \RegFile/_3595_ ;
wire \RegFile/_3596_ ;
wire \RegFile/_3597_ ;
wire \RegFile/_3598_ ;
wire \RegFile/_3599_ ;
wire \RegFile/_3600_ ;
wire \RegFile/_3601_ ;
wire \RegFile/_3602_ ;
wire \RegFile/_3603_ ;
wire \RegFile/_3604_ ;
wire \RegFile/_3605_ ;
wire \RegFile/_3606_ ;
wire \RegFile/_3607_ ;
wire \RegFile/_3608_ ;
wire \RegFile/_3609_ ;
wire \RegFile/_3610_ ;
wire \RegFile/_3611_ ;
wire \RegFile/_3612_ ;
wire \RegFile/_3613_ ;
wire \RegFile/_3614_ ;
wire \RegFile/_3615_ ;
wire \RegFile/_3616_ ;
wire \RegFile/_3617_ ;
wire \RegFile/_3618_ ;
wire \RegFile/_3619_ ;
wire \RegFile/_3620_ ;
wire \RegFile/_3621_ ;
wire \RegFile/_3622_ ;
wire \RegFile/_3623_ ;
wire \RegFile/_3624_ ;
wire \RegFile/_3625_ ;
wire \RegFile/_3626_ ;
wire \RegFile/_3627_ ;
wire \RegFile/_3628_ ;
wire \RegFile/_3629_ ;
wire \RegFile/_3630_ ;
wire \RegFile/_3631_ ;
wire \RegFile/_3632_ ;
wire \RegFile/_3633_ ;
wire \RegFile/_3634_ ;
wire \RegFile/_3635_ ;
wire \RegFile/_3636_ ;
wire \RegFile/_3637_ ;
wire \RegFile/_3638_ ;
wire \RegFile/_3639_ ;
wire \RegFile/_3640_ ;
wire \RegFile/_3641_ ;
wire \RegFile/_3642_ ;
wire \RegFile/_3643_ ;
wire \RegFile/_3644_ ;
wire \RegFile/_3645_ ;
wire \RegFile/_3646_ ;
wire \RegFile/_3647_ ;
wire \RegFile/_3648_ ;
wire \RegFile/_3649_ ;
wire \RegFile/_3650_ ;
wire \RegFile/_3651_ ;
wire \RegFile/_3652_ ;
wire \RegFile/_3653_ ;
wire \RegFile/_3654_ ;
wire \RegFile/_3655_ ;
wire \RegFile/_3656_ ;
wire \RegFile/_3657_ ;
wire \RegFile/_3658_ ;
wire \RegFile/_3659_ ;
wire \RegFile/_3660_ ;
wire \RegFile/_3661_ ;
wire \RegFile/_3662_ ;
wire \RegFile/_3663_ ;
wire \RegFile/_3664_ ;
wire \RegFile/_3665_ ;
wire \RegFile/_3666_ ;
wire \RegFile/_3667_ ;
wire \RegFile/_3668_ ;
wire \RegFile/_3669_ ;
wire \RegFile/_3670_ ;
wire \RegFile/_3671_ ;
wire \RegFile/_3672_ ;
wire \RegFile/_3673_ ;
wire \RegFile/_3674_ ;
wire \RegFile/_3675_ ;
wire \RegFile/_3676_ ;
wire \RegFile/_3677_ ;
wire \RegFile/_3678_ ;
wire \RegFile/_3679_ ;
wire \RegFile/_3680_ ;
wire \RegFile/_3681_ ;
wire \RegFile/_3682_ ;
wire \RegFile/_3683_ ;
wire \RegFile/_3684_ ;
wire \RegFile/_3685_ ;
wire \RegFile/_3686_ ;
wire \RegFile/_3687_ ;
wire \RegFile/_3688_ ;
wire \RegFile/_3689_ ;
wire \RegFile/_3690_ ;
wire \RegFile/_3691_ ;
wire \RegFile/_3692_ ;
wire \RegFile/_3693_ ;
wire \RegFile/_3694_ ;
wire \RegFile/_3695_ ;
wire \RegFile/_3696_ ;
wire \RegFile/_3697_ ;
wire \RegFile/_3698_ ;
wire \RegFile/_3699_ ;
wire \RegFile/_3700_ ;
wire \RegFile/_3701_ ;
wire \RegFile/_3702_ ;
wire \RegFile/_3703_ ;
wire \RegFile/_3704_ ;
wire \RegFile/_3705_ ;
wire \RegFile/_3706_ ;
wire \RegFile/_3707_ ;
wire \RegFile/_3708_ ;
wire \RegFile/_3709_ ;
wire \RegFile/_3710_ ;
wire \RegFile/_3711_ ;
wire \RegFile/_3712_ ;
wire \RegFile/_3713_ ;
wire \RegFile/_3714_ ;
wire \RegFile/_3715_ ;
wire \RegFile/_3716_ ;
wire \RegFile/_3717_ ;
wire \RegFile/_3718_ ;
wire \RegFile/_3719_ ;
wire \RegFile/_3720_ ;
wire \RegFile/_3721_ ;
wire \RegFile/_3722_ ;
wire \RegFile/_3723_ ;
wire \RegFile/_3724_ ;
wire \RegFile/_3725_ ;
wire \RegFile/_3726_ ;
wire \RegFile/_3727_ ;
wire \RegFile/_3728_ ;
wire \RegFile/_3729_ ;
wire \RegFile/_3730_ ;
wire \RegFile/_3731_ ;
wire \RegFile/_3732_ ;
wire \RegFile/_3733_ ;
wire \RegFile/_3734_ ;
wire \RegFile/_3735_ ;
wire \RegFile/_3736_ ;
wire \RegFile/_3737_ ;
wire \RegFile/_3738_ ;
wire \RegFile/_3739_ ;
wire \RegFile/_3740_ ;
wire \RegFile/_3741_ ;
wire \RegFile/_3742_ ;
wire \RegFile/_3743_ ;
wire \RegFile/_3744_ ;
wire \RegFile/_3745_ ;
wire \RegFile/_3746_ ;
wire \RegFile/_3747_ ;
wire \RegFile/_3748_ ;
wire \RegFile/_3749_ ;
wire \RegFile/_3750_ ;
wire \RegFile/_3751_ ;
wire \RegFile/_3752_ ;
wire \RegFile/_3753_ ;
wire \RegFile/_3754_ ;
wire \RegFile/_3755_ ;
wire \RegFile/_3756_ ;
wire \RegFile/_3757_ ;
wire \RegFile/_3758_ ;
wire \RegFile/_3759_ ;
wire \RegFile/_3760_ ;
wire \RegFile/_3761_ ;
wire \RegFile/_3762_ ;
wire \RegFile/_3763_ ;
wire \RegFile/_3764_ ;
wire \RegFile/_3765_ ;
wire \RegFile/_3766_ ;
wire \RegFile/_3767_ ;
wire \RegFile/_3768_ ;
wire \RegFile/_3769_ ;
wire \RegFile/_3770_ ;
wire \RegFile/_3771_ ;
wire \RegFile/_3772_ ;
wire \RegFile/_3773_ ;
wire \RegFile/_3774_ ;
wire \RegFile/_3775_ ;
wire \RegFile/_3776_ ;
wire \RegFile/_3777_ ;
wire \RegFile/_3778_ ;
wire \RegFile/_3779_ ;
wire \RegFile/_3780_ ;
wire \RegFile/_3781_ ;
wire \RegFile/_3782_ ;
wire \RegFile/_3783_ ;
wire \RegFile/_3784_ ;
wire \RegFile/_3785_ ;
wire \RegFile/_3786_ ;
wire \RegFile/_3787_ ;
wire \RegFile/_3788_ ;
wire \RegFile/_3789_ ;
wire \RegFile/_3790_ ;
wire \RegFile/_3791_ ;
wire \RegFile/_3792_ ;
wire \RegFile/_3793_ ;
wire \RegFile/_3794_ ;
wire \RegFile/_3795_ ;
wire \RegFile/_3796_ ;
wire \RegFile/_3797_ ;
wire \RegFile/_3798_ ;
wire \RegFile/_3799_ ;
wire \RegFile/_3800_ ;
wire \RegFile/_3801_ ;
wire \RegFile/_3802_ ;
wire \RegFile/_3803_ ;
wire \RegFile/_3804_ ;
wire \RegFile/_3805_ ;
wire \RegFile/_3806_ ;
wire \RegFile/_3807_ ;
wire \RegFile/_3808_ ;
wire \RegFile/_3809_ ;
wire \RegFile/_3810_ ;
wire \RegFile/_3811_ ;
wire \RegFile/_3812_ ;
wire \RegFile/_3813_ ;
wire \RegFile/_3814_ ;
wire \RegFile/_3815_ ;
wire \RegFile/_3816_ ;
wire \RegFile/_3817_ ;
wire \RegFile/_3818_ ;
wire \RegFile/_3819_ ;
wire \RegFile/_3820_ ;
wire \RegFile/_3821_ ;
wire \RegFile/_3822_ ;
wire \RegFile/_3823_ ;
wire \RegFile/_3824_ ;
wire \RegFile/_3825_ ;
wire \RegFile/_3826_ ;
wire \RegFile/_3827_ ;
wire \RegFile/_3828_ ;
wire \RegFile/_3829_ ;
wire \RegFile/_3830_ ;
wire \RegFile/_3831_ ;
wire \RegFile/_3832_ ;
wire \RegFile/_3833_ ;
wire \RegFile/_3834_ ;
wire \RegFile/_3835_ ;
wire \RegFile/_3836_ ;
wire \RegFile/_3837_ ;
wire \RegFile/_3838_ ;
wire \RegFile/_3839_ ;
wire \RegFile/_3840_ ;
wire \RegFile/_3841_ ;
wire \RegFile/_3842_ ;
wire \RegFile/_3843_ ;
wire \RegFile/_3844_ ;
wire \RegFile/_3845_ ;
wire \RegFile/_3846_ ;
wire \RegFile/_3847_ ;
wire \RegFile/_3848_ ;
wire \RegFile/_3849_ ;
wire \RegFile/_3850_ ;
wire \RegFile/_3851_ ;
wire \RegFile/_3852_ ;
wire \RegFile/_3853_ ;
wire \RegFile/_3854_ ;
wire \RegFile/_3855_ ;
wire \RegFile/_3856_ ;
wire \RegFile/_3857_ ;
wire \RegFile/_3858_ ;
wire \RegFile/_3859_ ;
wire \RegFile/_3860_ ;
wire \RegFile/_3861_ ;
wire \RegFile/_3862_ ;
wire \RegFile/_3863_ ;
wire \RegFile/_3864_ ;
wire \RegFile/_3865_ ;
wire \RegFile/_3866_ ;
wire \RegFile/_3867_ ;
wire \RegFile/_3868_ ;
wire \RegFile/_3869_ ;
wire \RegFile/_3870_ ;
wire \RegFile/_3871_ ;
wire \RegFile/_3872_ ;
wire \RegFile/_3873_ ;
wire \RegFile/_3874_ ;
wire \RegFile/_3875_ ;
wire \RegFile/_3876_ ;
wire \RegFile/_3877_ ;
wire \RegFile/_3878_ ;
wire \RegFile/_3879_ ;
wire \RegFile/_3880_ ;
wire \RegFile/_3881_ ;
wire \RegFile/_3882_ ;
wire \RegFile/_3883_ ;
wire \RegFile/_3884_ ;
wire \RegFile/_3885_ ;
wire \RegFile/_3886_ ;
wire \RegFile/_3887_ ;
wire \RegFile/_3888_ ;
wire \RegFile/_3889_ ;
wire \RegFile/_3890_ ;
wire \RegFile/_3891_ ;
wire \RegFile/_3892_ ;
wire \RegFile/_3893_ ;
wire \RegFile/_3894_ ;
wire \RegFile/_3895_ ;
wire \RegFile/_3896_ ;
wire \RegFile/_3897_ ;
wire \RegFile/_3898_ ;
wire \RegFile/_3899_ ;
wire \RegFile/_3900_ ;
wire \RegFile/_3901_ ;
wire \RegFile/_3902_ ;
wire \RegFile/_3903_ ;
wire \RegFile/_3904_ ;
wire \RegFile/_3905_ ;
wire \RegFile/_3906_ ;
wire \RegFile/_3907_ ;
wire \RegFile/_3908_ ;
wire \RegFile/_3909_ ;
wire \RegFile/_3910_ ;
wire \RegFile/_3911_ ;
wire \RegFile/_3912_ ;
wire \RegFile/_3913_ ;
wire \RegFile/_3914_ ;
wire \RegFile/_3915_ ;
wire \RegFile/_3916_ ;
wire \RegFile/_3917_ ;
wire \RegFile/_3918_ ;
wire \RegFile/_3919_ ;
wire \RegFile/_3920_ ;
wire \RegFile/_3921_ ;
wire \RegFile/_3922_ ;
wire \RegFile/_3923_ ;
wire \RegFile/_3924_ ;
wire \RegFile/_3925_ ;
wire \RegFile/_3926_ ;
wire \RegFile/_3927_ ;
wire \RegFile/_3928_ ;
wire \RegFile/_3929_ ;
wire \RegFile/_3930_ ;
wire \RegFile/_3931_ ;
wire \RegFile/_3932_ ;
wire \RegFile/_3933_ ;
wire \RegFile/_3934_ ;
wire \RegFile/_3935_ ;
wire \RegFile/_3936_ ;
wire \RegFile/_3937_ ;
wire \RegFile/_3938_ ;
wire \RegFile/_3939_ ;
wire \RegFile/_3940_ ;
wire \RegFile/_3941_ ;
wire \RegFile/_3942_ ;
wire \RegFile/_3943_ ;
wire \RegFile/_3944_ ;
wire \RegFile/_3945_ ;
wire \RegFile/_3946_ ;
wire \RegFile/_3947_ ;
wire \RegFile/_3948_ ;
wire \RegFile/_3949_ ;
wire \RegFile/_3950_ ;
wire \RegFile/_3951_ ;
wire \RegFile/_3952_ ;
wire \RegFile/_3953_ ;
wire \RegFile/_3954_ ;
wire \RegFile/_3955_ ;
wire \RegFile/_3956_ ;
wire \RegFile/_3957_ ;
wire \RegFile/_3958_ ;
wire \RegFile/_3959_ ;
wire \RegFile/_3960_ ;
wire \RegFile/_3961_ ;
wire \RegFile/_3962_ ;
wire \RegFile/_3963_ ;
wire \RegFile/_3964_ ;
wire \RegFile/_3965_ ;
wire \RegFile/_3966_ ;
wire \RegFile/_3967_ ;
wire \RegFile/_3968_ ;
wire \RegFile/_3969_ ;
wire \RegFile/_3970_ ;
wire \RegFile/_3971_ ;
wire \RegFile/_3972_ ;
wire \RegFile/_3973_ ;
wire \RegFile/_3974_ ;
wire \RegFile/_3975_ ;
wire \RegFile/_3976_ ;
wire \RegFile/_3977_ ;
wire \RegFile/_3978_ ;
wire \RegFile/_3979_ ;
wire \RegFile/_3980_ ;
wire \RegFile/_3981_ ;
wire \RegFile/_3982_ ;
wire \RegFile/_3983_ ;
wire \RegFile/_3984_ ;
wire \RegFile/_3985_ ;
wire \RegFile/_3986_ ;
wire \RegFile/_3987_ ;
wire \RegFile/_3988_ ;
wire \RegFile/_3989_ ;
wire \RegFile/_3990_ ;
wire \RegFile/_3991_ ;
wire \RegFile/_3992_ ;
wire \RegFile/_3993_ ;
wire \RegFile/_3994_ ;
wire \RegFile/_3995_ ;
wire \RegFile/_3996_ ;
wire \RegFile/_3997_ ;
wire \RegFile/_3998_ ;
wire \RegFile/_3999_ ;
wire \RegFile/_4000_ ;
wire \RegFile/_4001_ ;
wire \RegFile/_4002_ ;
wire \RegFile/_4003_ ;
wire \RegFile/_4004_ ;
wire \RegFile/_4005_ ;
wire \RegFile/_4006_ ;
wire \RegFile/_4007_ ;
wire \RegFile/_4008_ ;
wire \RegFile/_4009_ ;
wire \RegFile/_4010_ ;
wire \RegFile/_4011_ ;
wire \RegFile/_4012_ ;
wire \RegFile/_4013_ ;
wire \RegFile/_4014_ ;
wire \RegFile/_4015_ ;
wire \RegFile/_4016_ ;
wire \RegFile/_4017_ ;
wire \RegFile/_4018_ ;
wire \RegFile/_4019_ ;
wire \RegFile/_4020_ ;
wire \RegFile/_4021_ ;
wire \RegFile/_4022_ ;
wire \RegFile/_4023_ ;
wire \RegFile/_4024_ ;
wire \RegFile/_4025_ ;
wire \RegFile/_4026_ ;
wire \RegFile/_4027_ ;
wire \RegFile/_4028_ ;
wire \RegFile/_4029_ ;
wire \RegFile/_4030_ ;
wire \RegFile/_4031_ ;
wire \RegFile/_4032_ ;
wire \RegFile/_4033_ ;
wire \RegFile/_4034_ ;
wire \RegFile/_4035_ ;
wire \RegFile/_4036_ ;
wire \RegFile/_4037_ ;
wire \RegFile/_4038_ ;
wire \RegFile/_4039_ ;
wire \RegFile/_4040_ ;
wire \RegFile/_4041_ ;
wire \RegFile/_4042_ ;
wire \RegFile/_4043_ ;
wire \RegFile/_4044_ ;
wire \RegFile/_4045_ ;
wire \RegFile/_4046_ ;
wire \RegFile/_4047_ ;
wire \RegFile/_4048_ ;
wire \RegFile/_4049_ ;
wire \RegFile/_4050_ ;
wire \RegFile/_4051_ ;
wire \RegFile/_4052_ ;
wire \RegFile/_4053_ ;
wire \RegFile/_4054_ ;
wire \RegFile/_4055_ ;
wire \RegFile/_4056_ ;
wire \RegFile/_4057_ ;
wire \RegFile/_4058_ ;
wire \RegFile/_4059_ ;
wire \RegFile/_4060_ ;
wire \RegFile/_4061_ ;
wire \RegFile/_4062_ ;
wire \RegFile/_4063_ ;
wire \RegFile/_4064_ ;
wire \RegFile/_4065_ ;
wire \RegFile/_4066_ ;
wire \RegFile/_4067_ ;
wire \RegFile/_4068_ ;
wire \RegFile/_4069_ ;
wire \RegFile/_4070_ ;
wire \RegFile/_4071_ ;
wire \RegFile/_4072_ ;
wire \RegFile/_4073_ ;
wire \RegFile/_4074_ ;
wire \RegFile/_4075_ ;
wire \RegFile/_4076_ ;
wire \RegFile/_4077_ ;
wire \RegFile/_4078_ ;
wire \RegFile/_4079_ ;
wire \RegFile/_4080_ ;
wire \RegFile/_4081_ ;
wire \RegFile/_4082_ ;
wire \RegFile/_4083_ ;
wire \RegFile/_4084_ ;
wire \RegFile/_4085_ ;
wire \RegFile/_4086_ ;
wire \RegFile/_4087_ ;
wire \RegFile/_4088_ ;
wire \RegFile/_4089_ ;
wire \RegFile/_4090_ ;
wire \RegFile/_4091_ ;
wire \RegFile/_4092_ ;
wire \RegFile/_4093_ ;
wire \RegFile/_4094_ ;
wire \RegFile/_4095_ ;
wire \RegFile/_4096_ ;
wire \RegFile/_4097_ ;
wire \RegFile/_4098_ ;
wire \RegFile/_4099_ ;
wire \RegFile/_4100_ ;
wire \RegFile/_4101_ ;
wire \RegFile/_4102_ ;
wire \RegFile/_4103_ ;
wire \RegFile/_4104_ ;
wire \RegFile/_4105_ ;
wire \RegFile/_4106_ ;
wire \RegFile/_4107_ ;
wire \RegFile/_4108_ ;
wire \RegFile/_4109_ ;
wire \RegFile/_4110_ ;
wire \RegFile/_4111_ ;
wire \RegFile/_4112_ ;
wire \RegFile/_4113_ ;
wire \RegFile/_4114_ ;
wire \RegFile/_4115_ ;
wire \RegFile/_4116_ ;
wire \RegFile/_4117_ ;
wire \RegFile/_4118_ ;
wire \RegFile/_4119_ ;
wire \RegFile/_4120_ ;
wire \RegFile/_4121_ ;
wire \RegFile/_4122_ ;
wire \RegFile/_4123_ ;
wire \RegFile/_4124_ ;
wire \RegFile/_4125_ ;
wire \RegFile/_4126_ ;
wire \RegFile/_4127_ ;
wire \RegFile/_4128_ ;
wire \RegFile/_4129_ ;
wire \RegFile/_4130_ ;
wire \RegFile/_4131_ ;
wire \RegFile/_4132_ ;
wire \RegFile/_4133_ ;
wire \RegFile/_4134_ ;
wire \RegFile/_4135_ ;
wire \RegFile/_4136_ ;
wire \RegFile/_4137_ ;
wire \RegFile/_4138_ ;
wire \RegFile/_4139_ ;
wire \RegFile/_4140_ ;
wire \RegFile/_4141_ ;
wire \RegFile/_4142_ ;
wire \RegFile/_4143_ ;
wire \RegFile/_4144_ ;
wire \RegFile/_4145_ ;
wire \RegFile/_4146_ ;
wire \RegFile/_4147_ ;
wire \RegFile/_4148_ ;
wire \RegFile/_4149_ ;
wire \RegFile/_4150_ ;
wire \RegFile/_4151_ ;
wire \RegFile/_4152_ ;
wire \RegFile/_4153_ ;
wire \RegFile/_4154_ ;
wire \RegFile/_4155_ ;
wire \RegFile/_4156_ ;
wire \RegFile/_4157_ ;
wire \RegFile/_4158_ ;
wire \RegFile/_4159_ ;
wire \RegFile/_4160_ ;
wire \RegFile/_4161_ ;
wire \RegFile/_4162_ ;
wire \RegFile/_4163_ ;
wire \RegFile/_4164_ ;
wire \RegFile/_4165_ ;
wire \RegFile/_4166_ ;
wire \RegFile/_4167_ ;
wire \RegFile/_4168_ ;
wire \RegFile/_4169_ ;
wire \RegFile/_4170_ ;
wire \RegFile/_4171_ ;
wire \RegFile/_4172_ ;
wire \RegFile/_4173_ ;
wire \RegFile/_4174_ ;
wire \RegFile/_4175_ ;
wire \RegFile/_4176_ ;
wire \RegFile/_4177_ ;
wire \RegFile/_4178_ ;
wire \RegFile/_4179_ ;
wire \RegFile/_4180_ ;
wire \RegFile/_4181_ ;
wire \RegFile/_4182_ ;
wire \RegFile/_4183_ ;
wire \RegFile/_4184_ ;
wire \RegFile/_4185_ ;
wire \RegFile/_4186_ ;
wire \RegFile/_4187_ ;
wire \RegFile/_4188_ ;
wire \RegFile/_4189_ ;
wire \RegFile/_4190_ ;
wire \RegFile/_4191_ ;
wire \RegFile/_4192_ ;
wire \RegFile/_4193_ ;
wire \RegFile/_4194_ ;
wire \RegFile/_4195_ ;
wire \RegFile/_4196_ ;
wire \RegFile/_4197_ ;
wire \RegFile/_4198_ ;
wire \RegFile/_4199_ ;
wire \RegFile/_4200_ ;
wire \RegFile/_4201_ ;
wire \RegFile/_4202_ ;
wire \RegFile/_4203_ ;
wire \RegFile/_4204_ ;
wire \RegFile/_4205_ ;
wire \RegFile/_4206_ ;
wire \RegFile/_4207_ ;
wire \RegFile/_4208_ ;
wire \RegFile/_4209_ ;
wire \RegFile/_4210_ ;
wire \RegFile/_4211_ ;
wire \RegFile/_4212_ ;
wire \RegFile/_4213_ ;
wire \RegFile/_4214_ ;
wire \RegFile/_4215_ ;
wire \RegFile/_4216_ ;
wire \RegFile/_4217_ ;
wire \RegFile/_4218_ ;
wire \RegFile/_4219_ ;
wire \RegFile/_4220_ ;
wire \RegFile/_4221_ ;
wire \RegFile/_4222_ ;
wire \RegFile/_4223_ ;
wire \RegFile/_4224_ ;
wire \RegFile/_4225_ ;
wire \RegFile/_4226_ ;
wire \RegFile/_4227_ ;
wire \RegFile/_4228_ ;
wire \RegFile/_4229_ ;
wire \RegFile/_4230_ ;
wire \RegFile/_4231_ ;
wire \RegFile/_4232_ ;
wire \RegFile/_4233_ ;
wire \RegFile/_4234_ ;
wire \RegFile/_4235_ ;
wire \RegFile/_4236_ ;
wire \RegFile/_4237_ ;
wire \RegFile/_4238_ ;
wire \RegFile/_4239_ ;
wire \RegFile/_4240_ ;
wire \RegFile/_4241_ ;
wire \RegFile/_4242_ ;
wire \RegFile/_4243_ ;
wire \RegFile/_4244_ ;
wire \RegFile/_4245_ ;
wire \RegFile/_4246_ ;
wire \RegFile/_4247_ ;
wire \RegFile/_4248_ ;
wire \RegFile/_4249_ ;
wire \RegFile/_4250_ ;
wire \RegFile/_4251_ ;
wire \RegFile/_4252_ ;
wire \RegFile/_4253_ ;
wire \RegFile/_4254_ ;
wire \RegFile/_4255_ ;
wire \RegFile/_4256_ ;
wire \RegFile/_4257_ ;
wire \RegFile/_4258_ ;
wire \RegFile/_4259_ ;
wire \RegFile/_4260_ ;
wire \RegFile/_4261_ ;
wire \RegFile/_4262_ ;
wire \RegFile/_4263_ ;
wire \RegFile/_4264_ ;
wire \RegFile/_4265_ ;
wire \RegFile/_4266_ ;
wire \RegFile/_4267_ ;
wire \RegFile/_4268_ ;
wire \RegFile/_4269_ ;
wire \RegFile/_4270_ ;
wire \RegFile/_4271_ ;
wire \RegFile/_4272_ ;
wire \RegFile/_4273_ ;
wire \RegFile/_4274_ ;
wire \RegFile/_4275_ ;
wire \RegFile/_4276_ ;
wire \RegFile/_4277_ ;
wire \RegFile/_4278_ ;
wire \RegFile/_4279_ ;
wire \RegFile/_4280_ ;
wire \RegFile/_4281_ ;
wire \RegFile/_4282_ ;
wire \RegFile/_4283_ ;
wire \RegFile/_4284_ ;
wire \RegFile/_4285_ ;
wire \RegFile/_4286_ ;
wire \RegFile/_4287_ ;
wire \RegFile/_4288_ ;
wire \RegFile/_4289_ ;
wire \RegFile/_4290_ ;
wire \RegFile/_4291_ ;
wire \RegFile/_4292_ ;
wire \RegFile/_4293_ ;
wire \RegFile/_4294_ ;
wire \RegFile/_4295_ ;
wire \RegFile/_4296_ ;
wire \RegFile/_4297_ ;
wire \RegFile/_4298_ ;
wire \RegFile/_4299_ ;
wire \RegFile/_4300_ ;
wire \RegFile/_4301_ ;
wire \RegFile/_4302_ ;
wire \RegFile/_4303_ ;
wire \RegFile/_4304_ ;
wire \RegFile/_4305_ ;
wire \RegFile/_4306_ ;
wire \RegFile/_4307_ ;
wire \RegFile/_4308_ ;
wire \RegFile/_4309_ ;
wire \RegFile/_4310_ ;
wire \RegFile/_4311_ ;
wire \RegFile/_4312_ ;
wire \RegFile/_4313_ ;
wire \RegFile/_4314_ ;
wire \RegFile/_4315_ ;
wire \RegFile/_4316_ ;
wire \RegFile/_4317_ ;
wire \RegFile/_4318_ ;
wire \RegFile/_4319_ ;
wire \RegFile/_4320_ ;
wire \RegFile/_4321_ ;
wire \RegFile/_4322_ ;
wire \RegFile/_4323_ ;
wire \RegFile/_4324_ ;
wire \RegFile/_4325_ ;
wire \RegFile/_4326_ ;
wire \RegFile/_4327_ ;
wire \RegFile/_4328_ ;
wire \RegFile/_4329_ ;
wire \RegFile/_4330_ ;
wire \RegFile/_4331_ ;
wire \RegFile/_4332_ ;
wire \RegFile/_4333_ ;
wire \RegFile/_4334_ ;
wire \RegFile/_4335_ ;
wire \RegFile/_4336_ ;
wire \RegFile/_4337_ ;
wire \RegFile/_4338_ ;
wire \RegFile/_4339_ ;
wire \RegFile/_4340_ ;
wire \RegFile/_4341_ ;
wire \RegFile/_4342_ ;
wire \RegFile/_4343_ ;
wire \RegFile/_4344_ ;
wire \RegFile/_4345_ ;
wire \RegFile/_4346_ ;
wire \RegFile/_4347_ ;
wire \RegFile/_4348_ ;
wire \RegFile/_4349_ ;
wire \RegFile/_4350_ ;
wire \RegFile/_4351_ ;
wire \RegFile/_4352_ ;
wire \RegFile/_4353_ ;
wire \RegFile/_4354_ ;
wire \RegFile/_4355_ ;
wire \RegFile/_4356_ ;
wire \RegFile/_4357_ ;
wire \RegFile/_4358_ ;
wire \RegFile/_4359_ ;
wire \RegFile/_4360_ ;
wire \RegFile/_4361_ ;
wire \RegFile/_4362_ ;
wire \RegFile/_4363_ ;
wire \RegFile/_4364_ ;
wire \RegFile/_4365_ ;
wire \RegFile/_4366_ ;
wire \RegFile/_4367_ ;
wire \RegFile/_4368_ ;
wire \RegFile/_4369_ ;
wire \RegFile/_4370_ ;
wire \RegFile/_4371_ ;
wire \RegFile/_4372_ ;
wire \RegFile/_4373_ ;
wire \RegFile/_4374_ ;
wire \RegFile/_4375_ ;
wire \RegFile/_4376_ ;
wire \RegFile/_4377_ ;
wire \RegFile/_4378_ ;
wire \RegFile/_4379_ ;
wire \RegFile/_4380_ ;
wire \RegFile/_4381_ ;
wire \RegFile/_4382_ ;
wire \RegFile/_4383_ ;
wire \RegFile/_4384_ ;
wire \RegFile/_4385_ ;
wire \RegFile/_4386_ ;
wire \RegFile/_4387_ ;
wire \RegFile/_4388_ ;
wire \RegFile/_4389_ ;
wire \RegFile/_4390_ ;
wire \RegFile/_4391_ ;
wire \RegFile/_4392_ ;
wire \RegFile/_4393_ ;
wire \RegFile/_4394_ ;
wire \RegFile/_4395_ ;
wire \RegFile/_4396_ ;
wire \RegFile/_4397_ ;
wire \RegFile/_4398_ ;
wire \RegFile/_4399_ ;
wire \RegFile/_4400_ ;
wire \RegFile/_4401_ ;
wire \RegFile/_4402_ ;
wire \RegFile/_4403_ ;
wire \RegFile/_4404_ ;
wire \RegFile/_4405_ ;
wire \RegFile/_4406_ ;
wire \RegFile/_4407_ ;
wire \RegFile/_4408_ ;
wire \RegFile/_4409_ ;
wire \RegFile/_4410_ ;
wire \RegFile/_4411_ ;
wire \RegFile/_4412_ ;
wire \RegFile/_4413_ ;
wire \RegFile/_4414_ ;
wire \RegFile/_4415_ ;
wire \RegFile/_4416_ ;
wire \RegFile/_4417_ ;
wire \RegFile/_4418_ ;
wire \RegFile/_4419_ ;
wire \RegFile/_4420_ ;
wire \RegFile/_4421_ ;
wire \RegFile/_4422_ ;
wire \RegFile/_4423_ ;
wire \RegFile/_4424_ ;
wire \RegFile/_4425_ ;
wire \RegFile/_4426_ ;
wire \RegFile/_4427_ ;
wire \RegFile/_4428_ ;
wire \RegFile/_4429_ ;
wire \RegFile/_4430_ ;
wire \RegFile/_4431_ ;
wire \RegFile/_4432_ ;
wire \RegFile/_4433_ ;
wire \RegFile/_4434_ ;
wire \RegFile/_4435_ ;
wire \RegFile/_4436_ ;
wire \RegFile/_4437_ ;
wire \RegFile/_4438_ ;
wire \RegFile/_4439_ ;
wire \RegFile/_4440_ ;
wire \RegFile/_4441_ ;
wire \RegFile/_4442_ ;
wire \RegFile/_4443_ ;
wire \RegFile/_4444_ ;
wire \RegFile/_4445_ ;
wire \RegFile/_4446_ ;
wire \RegFile/_4447_ ;
wire \RegFile/_4448_ ;
wire \RegFile/_4449_ ;
wire \RegFile/_4450_ ;
wire \RegFile/_4451_ ;
wire \RegFile/_4452_ ;
wire \RegFile/_4453_ ;
wire \RegFile/_4454_ ;
wire \RegFile/_4455_ ;
wire \RegFile/_4456_ ;
wire \RegFile/_4457_ ;
wire \RegFile/_4458_ ;
wire \RegFile/_4459_ ;
wire \RegFile/_4460_ ;
wire \RegFile/_4461_ ;
wire \RegFile/_4462_ ;
wire \RegFile/_4463_ ;
wire \RegFile/_4464_ ;
wire \RegFile/_4465_ ;
wire \RegFile/_4466_ ;
wire \RegFile/_4467_ ;
wire \RegFile/_4468_ ;
wire \RegFile/_4469_ ;
wire \RegFile/_4470_ ;
wire \RegFile/_4471_ ;
wire \RegFile/_4472_ ;
wire \RegFile/_4473_ ;
wire \RegFile/_4474_ ;
wire \RegFile/_4475_ ;
wire \RegFile/_4476_ ;
wire \RegFile/_4477_ ;
wire \RegFile/_4478_ ;
wire \RegFile/_4479_ ;
wire \RegFile/_4480_ ;
wire \RegFile/_4481_ ;
wire \RegFile/_4482_ ;
wire \RegFile/_4483_ ;
wire \RegFile/_4484_ ;
wire \RegFile/_4485_ ;
wire \RegFile/_4486_ ;
wire \RegFile/_4487_ ;
wire \RegFile/_4488_ ;
wire \RegFile/_4489_ ;
wire \RegFile/_4490_ ;
wire \RegFile/_4491_ ;
wire \RegFile/_4492_ ;
wire \RegFile/_4493_ ;
wire \RegFile/_4494_ ;
wire \RegFile/_4495_ ;
wire \RegFile/_4496_ ;
wire \RegFile/_4497_ ;
wire \RegFile/_4498_ ;
wire \RegFile/_4499_ ;
wire \RegFile/_4500_ ;
wire \RegFile/_4501_ ;
wire \RegFile/_4502_ ;
wire \RegFile/_4503_ ;
wire \RegFile/_4504_ ;
wire \RegFile/_4505_ ;
wire \RegFile/_4506_ ;
wire \RegFile/_4507_ ;
wire \RegFile/_4508_ ;
wire \RegFile/_4509_ ;
wire \RegFile/_4510_ ;
wire \RegFile/_4511_ ;
wire \RegFile/_4512_ ;
wire \RegFile/_4513_ ;
wire \RegFile/_4514_ ;
wire \RegFile/_4515_ ;
wire \RegFile/_4516_ ;
wire \RegFile/_4517_ ;
wire \RegFile/_4518_ ;
wire \RegFile/_4519_ ;
wire \RegFile/_4520_ ;
wire \RegFile/_4521_ ;
wire \RegFile/_4522_ ;
wire \RegFile/_4523_ ;
wire \RegFile/_4524_ ;
wire \RegFile/_4525_ ;
wire \RegFile/_4526_ ;
wire \RegFile/_4527_ ;
wire \RegFile/_4528_ ;
wire \RegFile/_4529_ ;
wire \RegFile/_4530_ ;
wire \RegFile/_4531_ ;
wire \RegFile/_4532_ ;
wire \RegFile/_4533_ ;
wire \RegFile/_4534_ ;
wire \RegFile/_4535_ ;
wire \RegFile/_4536_ ;
wire \RegFile/_4537_ ;
wire \RegFile/_4538_ ;
wire \RegFile/_4539_ ;
wire \RegFile/_4540_ ;
wire \RegFile/_4541_ ;
wire \RegFile/_4542_ ;
wire \RegFile/_4543_ ;
wire \RegFile/_4544_ ;
wire \RegFile/_4545_ ;
wire \RegFile/_4546_ ;
wire \RegFile/_4547_ ;
wire \RegFile/_4548_ ;
wire \RegFile/_4549_ ;
wire \RegFile/_4550_ ;
wire \RegFile/_4551_ ;
wire \RegFile/_4552_ ;
wire \RegFile/_4553_ ;
wire \RegFile/_4554_ ;
wire \RegFile/_4555_ ;
wire \RegFile/_4556_ ;
wire \RegFile/_4557_ ;
wire \RegFile/_4558_ ;
wire \RegFile/_4559_ ;
wire \RegFile/_4560_ ;
wire \RegFile/_4561_ ;
wire \RegFile/_4562_ ;
wire \RegFile/_4563_ ;
wire \RegFile/_4564_ ;
wire \RegFile/_4565_ ;
wire \RegFile/_4566_ ;
wire \RegFile/_4567_ ;
wire \RegFile/_4568_ ;
wire \RegFile/_4569_ ;
wire \RegFile/_4570_ ;
wire \RegFile/_4571_ ;
wire \RegFile/_4572_ ;
wire \RegFile/_4573_ ;
wire \RegFile/_4574_ ;
wire \RegFile/_4575_ ;
wire \RegFile/_4576_ ;
wire \RegFile/_4577_ ;
wire \RegFile/_4578_ ;
wire \RegFile/_4579_ ;
wire \RegFile/_4580_ ;
wire \RegFile/_4581_ ;
wire \RegFile/_4582_ ;
wire \RegFile/_4583_ ;
wire \RegFile/_4584_ ;
wire \RegFile/_4585_ ;
wire \RegFile/_4586_ ;
wire \RegFile/_4587_ ;
wire \RegFile/_4588_ ;
wire \RegFile/_4589_ ;
wire \RegFile/_4590_ ;
wire \RegFile/_4591_ ;
wire \RegFile/_4592_ ;
wire \RegFile/_4593_ ;
wire \RegFile/_4594_ ;
wire \RegFile/_4595_ ;
wire \RegFile/_4596_ ;
wire \RegFile/_4597_ ;
wire \RegFile/_4598_ ;
wire \RegFile/_4599_ ;
wire \RegFile/_4600_ ;
wire \RegFile/_4601_ ;
wire \RegFile/_4602_ ;
wire \RegFile/_4603_ ;
wire \RegFile/_4604_ ;
wire \RegFile/_4605_ ;
wire \RegFile/_4606_ ;
wire \RegFile/_4607_ ;
wire \RegFile/_4608_ ;
wire \RegFile/_4609_ ;
wire \RegFile/_4610_ ;
wire \RegFile/_4611_ ;
wire \RegFile/_4612_ ;
wire \RegFile/_4613_ ;
wire \RegFile/_4614_ ;
wire \RegFile/_4615_ ;
wire \RegFile/_4616_ ;
wire \RegFile/_4617_ ;
wire \RegFile/_4618_ ;
wire \RegFile/_4619_ ;
wire \RegFile/_4620_ ;
wire \RegFile/_4621_ ;
wire \RegFile/_4622_ ;
wire \RegFile/_4623_ ;
wire \RegFile/_4624_ ;
wire \RegFile/_4625_ ;
wire \RegFile/_4626_ ;
wire \RegFile/_4627_ ;
wire \RegFile/_4628_ ;
wire \RegFile/_4629_ ;
wire \RegFile/_4630_ ;
wire \RegFile/_4631_ ;
wire \RegFile/_4632_ ;
wire \RegFile/_4633_ ;
wire \RegFile/_4634_ ;
wire \RegFile/_4635_ ;
wire \RegFile/_4636_ ;
wire \RegFile/_4637_ ;
wire \RegFile/_4638_ ;
wire \RegFile/_4639_ ;
wire \RegFile/_4640_ ;
wire \RegFile/_4641_ ;
wire \RegFile/_4642_ ;
wire \RegFile/_4643_ ;
wire \RegFile/_4644_ ;
wire \RegFile/_4645_ ;
wire \RegFile/_4646_ ;
wire \RegFile/_4647_ ;
wire \RegFile/_4648_ ;
wire \RegFile/_4649_ ;
wire \RegFile/_4650_ ;
wire \RegFile/_4651_ ;
wire \RegFile/_4652_ ;
wire \RegFile/_4653_ ;
wire \RegFile/_4654_ ;
wire \RegFile/_4655_ ;
wire \RegFile/_4656_ ;
wire \RegFile/_4657_ ;
wire \RegFile/_4658_ ;
wire \RegFile/_4659_ ;
wire \RegFile/_4660_ ;
wire \RegFile/_4661_ ;
wire \RegFile/_4662_ ;
wire \RegFile/_4663_ ;
wire \RegFile/_4664_ ;
wire \RegFile/_4665_ ;
wire \RegFile/_4666_ ;
wire \RegFile/_4667_ ;
wire \RegFile/_4668_ ;
wire \RegFile/_4669_ ;
wire \RegFile/_4670_ ;
wire \RegFile/_4671_ ;
wire \RegFile/_4672_ ;
wire \RegFile/_4673_ ;
wire \RegFile/_4674_ ;
wire \RegFile/_4675_ ;
wire \RegFile/_4676_ ;
wire \RegFile/_4677_ ;
wire \RegFile/_4678_ ;
wire \RegFile/_4679_ ;
wire \RegFile/_4680_ ;
wire \RegFile/_4681_ ;
wire \RegFile/_4682_ ;
wire \RegFile/_4683_ ;
wire \RegFile/_4684_ ;
wire \RegFile/_4685_ ;
wire \RegFile/_4686_ ;
wire \RegFile/_4687_ ;
wire \RegFile/_4688_ ;
wire \RegFile/_4689_ ;
wire \RegFile/_4690_ ;
wire \RegFile/_4691_ ;
wire \RegFile/_4692_ ;
wire \RegFile/_4693_ ;
wire \RegFile/_4694_ ;
wire \RegFile/_4695_ ;
wire \RegFile/_4696_ ;
wire \RegFile/_4697_ ;
wire \RegFile/_4698_ ;
wire \RegFile/_4699_ ;
wire \RegFile/_4700_ ;
wire \RegFile/_4701_ ;
wire \RegFile/_4702_ ;
wire \RegFile/_4703_ ;
wire \RegFile/_4704_ ;
wire \RegFile/_4705_ ;
wire \RegFile/_4706_ ;
wire \RegFile/_4707_ ;
wire \RegFile/_4708_ ;
wire \RegFile/_4709_ ;
wire \RegFile/_4710_ ;
wire \RegFile/_4711_ ;
wire \RegFile/_4712_ ;
wire \RegFile/_4713_ ;
wire \RegFile/_4714_ ;
wire \RegFile/_4715_ ;
wire \RegFile/_4716_ ;
wire \RegFile/_4717_ ;
wire \RegFile/_4718_ ;
wire \RegFile/_4719_ ;
wire \RegFile/_4720_ ;
wire \RegFile/_4721_ ;
wire \RegFile/_4722_ ;
wire \RegFile/_4723_ ;
wire \RegFile/_4724_ ;
wire \RegFile/_4725_ ;
wire \RegFile/_4726_ ;
wire \RegFile/_4727_ ;
wire \RegFile/_4728_ ;
wire \RegFile/_4729_ ;
wire \RegFile/_4730_ ;
wire \RegFile/_4731_ ;
wire \RegFile/_4732_ ;
wire \RegFile/_4733_ ;
wire \RegFile/_4734_ ;
wire \RegFile/_4735_ ;
wire \RegFile/_4736_ ;
wire \RegFile/_4737_ ;
wire \RegFile/_4738_ ;
wire \RegFile/_4739_ ;
wire \RegFile/_4740_ ;
wire \RegFile/_4741_ ;
wire \RegFile/_4742_ ;
wire \RegFile/_4743_ ;
wire \RegFile/_4744_ ;
wire \RegFile/_4745_ ;
wire \RegFile/_4746_ ;
wire \RegFile/_4747_ ;
wire \RegFile/_4748_ ;
wire \RegFile/_4749_ ;
wire \RegFile/_4750_ ;
wire \RegFile/_4751_ ;
wire \RegFile/_4752_ ;
wire \RegFile/_4753_ ;
wire \WBU/_000_ ;
wire \WBU/_001_ ;
wire \WBU/_002_ ;
wire \WBU/_003_ ;
wire \WBU/_004_ ;
wire \WBU/_005_ ;
wire \WBU/_006_ ;
wire \WBU/_007_ ;
wire \WBU/_008_ ;
wire \WBU/_009_ ;
wire \WBU/_010_ ;
wire \WBU/_011_ ;
wire \WBU/_012_ ;
wire \WBU/_013_ ;
wire \WBU/_014_ ;
wire \WBU/_015_ ;
wire \WBU/_016_ ;
wire \WBU/_017_ ;
wire \WBU/_018_ ;
wire \WBU/_019_ ;
wire \WBU/_020_ ;
wire \WBU/_021_ ;
wire \WBU/_022_ ;
wire \WBU/_023_ ;
wire \WBU/_024_ ;
wire \WBU/_025_ ;
wire \WBU/_026_ ;
wire \WBU/_027_ ;
wire \WBU/_028_ ;
wire \WBU/_029_ ;
wire \WBU/_030_ ;
wire \WBU/_031_ ;
wire \WBU/_032_ ;
wire \WBU/_033_ ;
wire \WBU/_034_ ;
wire \WBU/_035_ ;
wire \WBU/_036_ ;
wire \WBU/_037_ ;
wire \WBU/_038_ ;
wire \WBU/_039_ ;
wire \WBU/_040_ ;
wire \WBU/_041_ ;
wire \WBU/_042_ ;
wire \WBU/_043_ ;
wire \WBU/_044_ ;
wire \WBU/_045_ ;
wire \WBU/_046_ ;
wire \WBU/_047_ ;
wire \WBU/_048_ ;
wire \WBU/_049_ ;
wire \WBU/_050_ ;
wire \WBU/_051_ ;
wire \WBU/_052_ ;
wire \WBU/_053_ ;
wire \WBU/_054_ ;
wire \WBU/_055_ ;
wire \WBU/_056_ ;
wire \WBU/_057_ ;
wire \WBU/_058_ ;
wire \WBU/_059_ ;
wire \WBU/_060_ ;
wire \WBU/_061_ ;
wire \WBU/_062_ ;
wire \WBU/_063_ ;
wire \WBU/_064_ ;
wire \WBU/_065_ ;
wire \WBU/_066_ ;
wire \WBU/_067_ ;
wire \WBU/_068_ ;
wire \WBU/_069_ ;
wire \WBU/_070_ ;
wire \WBU/_071_ ;
wire \WBU/_072_ ;
wire \WBU/_073_ ;
wire \WBU/_074_ ;
wire \WBU/_075_ ;
wire \WBU/_076_ ;
wire \WBU/_077_ ;
wire \WBU/_078_ ;
wire \WBU/_079_ ;
wire \WBU/_080_ ;
wire \WBU/_081_ ;
wire \WBU/_082_ ;
wire \WBU/_083_ ;
wire \WBU/_084_ ;
wire \WBU/_085_ ;
wire \WBU/_086_ ;
wire \WBU/_087_ ;
wire \WBU/_088_ ;
wire \WBU/_089_ ;
wire \WBU/_090_ ;
wire \WBU/_091_ ;
wire \WBU/_092_ ;
wire \WBU/_093_ ;
wire \WBU/_094_ ;
wire \WBU/_095_ ;
wire \WBU/_096_ ;
wire \WBU/_097_ ;
wire \WBU/_098_ ;
wire \WBU/_099_ ;
wire \WBU/_100_ ;
wire \WBU/_101_ ;
wire \WBU/_102_ ;
wire \WBU/_103_ ;
wire \WBU/_104_ ;
wire \WBU/_105_ ;
wire \WBU/_106_ ;
wire \WBU/_107_ ;
wire \WBU/_108_ ;
wire \WBU/_109_ ;
wire \WBU/_110_ ;
wire \WBU/_111_ ;
wire \WBU/_112_ ;
wire \WBU/_113_ ;
wire \WBU/_114_ ;
wire \WBU/_115_ ;
wire \WBU/_116_ ;
wire \WBU/_117_ ;
wire \WBU/_118_ ;
wire \WBU/_119_ ;
wire \WBU/_120_ ;
wire \WBU/_121_ ;
wire \WBU/_122_ ;
wire \WBU/_123_ ;
wire \WBU/_124_ ;
wire \WBU/_125_ ;
wire \WBU/_126_ ;
wire \WBU/_127_ ;
wire \WBU/_128_ ;
wire \WBU/_129_ ;
wire \WBU/_130_ ;
wire \WBU/_131_ ;
wire \WBU/_132_ ;
wire \WBU/_133_ ;
wire \WBU/_134_ ;
wire \WBU/_135_ ;
wire \WBU/_136_ ;
wire \WBU/_137_ ;
wire \WBU/_138_ ;
wire \WBU/_139_ ;
wire \WBU/_140_ ;
wire \WBU/_141_ ;
wire \WBU/_142_ ;
wire \WBU/_143_ ;
wire \WBU/_144_ ;
wire \WBU/_145_ ;
wire \WBU/_146_ ;
wire \WBU/_147_ ;
wire \WBU/_148_ ;
wire \WBU/_149_ ;
wire \WBU/_150_ ;
wire \WBU/_151_ ;
wire \WBU/_152_ ;
wire \WBU/_153_ ;
wire \WBU/_154_ ;
wire \WBU/_155_ ;
wire \WBU/_156_ ;
wire \WBU/_157_ ;
wire \WBU/_158_ ;
wire \WBU/_159_ ;
wire \WBU/_160_ ;
wire \WBU/_161_ ;
wire \WBU/_162_ ;
wire \WBU/_163_ ;
wire \WBU/_164_ ;
wire \WBU/_165_ ;
wire \WBU/_166_ ;
wire \WBU/_167_ ;
wire \WBU/_168_ ;
wire \WBU/_169_ ;
wire \WBU/_170_ ;
wire \WBU/_171_ ;
wire \WBU/_172_ ;
wire \WBU/_173_ ;
wire \WBU/_174_ ;
wire \WBU/_175_ ;
wire \WBU/_176_ ;
wire \WBU/_177_ ;
wire \WBU/_178_ ;
wire \WBU/_179_ ;
wire \WBU/_180_ ;
wire \WBU/_181_ ;
wire \WBU/_182_ ;
wire \WBU/_183_ ;
wire \WBU/_184_ ;
wire \WBU/_185_ ;
wire \WBU/_186_ ;
wire \WBU/_187_ ;
wire \WBU/_188_ ;
wire \WBU/_189_ ;
wire \WBU/_190_ ;
wire \WBU/_191_ ;
wire \WBU/_192_ ;
wire \WBU/_193_ ;
wire \WBU/_194_ ;
wire \WBU/_195_ ;
wire \WBU/_196_ ;
wire \WBU/_197_ ;
wire \WBU/_198_ ;
wire \WBU/_199_ ;
wire \WBU/_200_ ;
wire \WBU/_201_ ;
wire \WBU/_202_ ;
wire \WBU/_203_ ;
wire \WBU/_204_ ;
wire \WBU/_205_ ;
wire \WBU/_206_ ;
wire \WBU/_207_ ;
wire \WBU/_208_ ;
wire \WBU/_209_ ;
wire \WBU/_210_ ;
wire \WBU/_211_ ;
wire \WBU/_212_ ;
wire \WBU/_213_ ;
wire \WBU/_214_ ;
wire \WBU/_215_ ;
wire \WBU/_216_ ;
wire \WBU/_217_ ;
wire \WBU/_218_ ;
wire \WBU/_219_ ;
wire \WBU/_220_ ;
wire \WBU/_221_ ;
wire \WBU/_222_ ;
wire \WBU/_223_ ;
wire \WBU/_224_ ;
wire \WBU/_225_ ;
wire \WBU/_226_ ;
wire \WBU/_227_ ;
wire \WBU/_228_ ;
wire \WBU/_229_ ;
wire \WBU/_230_ ;
wire \WBU/_231_ ;
wire \WBU/_232_ ;
wire \WBU/_233_ ;
wire \WBU/_234_ ;
wire \WBU/_235_ ;
wire \WBU/_236_ ;
wire \WBU/_237_ ;
wire \WBU/_238_ ;
wire \WBU/_239_ ;
wire \WBU/_240_ ;
wire \WBU/_241_ ;
wire \WBU/_242_ ;
wire \WBU/_243_ ;
wire \WBU/_244_ ;
wire \WBU/_245_ ;
wire \WBU/_246_ ;
wire \WBU/_247_ ;
wire \WBU/_248_ ;
wire \WBU/_249_ ;
wire \WBU/_250_ ;
wire \WBU/_251_ ;
wire \WBU/_252_ ;
wire \WBU/_253_ ;
wire \WBU/_254_ ;
wire \WBU/_255_ ;
wire \WBU/_256_ ;
wire \WBU/_257_ ;
wire \WBU/_258_ ;
wire \WBU/_259_ ;
wire \WBU/_260_ ;
wire \WBU/_261_ ;
wire \WBU/_262_ ;
wire \WBU/_263_ ;
wire \WBU/_264_ ;
wire \WBU/_265_ ;
wire \WBU/_266_ ;
wire \WBU/_267_ ;
wire \WBU/_268_ ;
wire \WBU/_269_ ;
wire \WBU/_270_ ;
wire \WBU/_271_ ;
wire \WBU/_272_ ;
wire \WBU/_273_ ;
wire \WBU/_274_ ;
wire fanout_net_1 ;
wire fanout_net_2 ;
wire fanout_net_3 ;
wire fanout_net_4 ;
wire fanout_net_5 ;
wire fanout_net_6 ;
wire fanout_net_7 ;
wire fanout_net_8 ;
wire fanout_net_9 ;
wire fanout_net_10 ;
wire fanout_net_11 ;
wire fanout_net_12 ;
wire fanout_net_13 ;
wire fanout_net_14 ;
wire fanout_net_15 ;
wire fanout_net_16 ;
wire fanout_net_17 ;
wire fanout_net_18 ;
wire fanout_net_19 ;
wire fanout_net_20 ;
wire [31:0] _AXI4Interconnect_io_fanIn_0_rdata ;
wire [1:0] _AXI4Interconnect_io_fanIn_0_rresp ;
wire [1:0] _AXI4Interconnect_io_fanIn_1_bresp ;
wire [31:0] _AXI4Interconnect_io_fanIn_1_rdata ;
wire [1:0] _AXI4Interconnect_io_fanIn_1_rresp ;
wire [31:0] _AXI4Interconnect_io_fanOut_0_araddr ;
wire [31:0] _AXI4Interconnect_io_fanOut_0_awaddr ;
wire [31:0] _AXI4Interconnect_io_fanOut_0_wdata ;
wire [1:0] _CLINT_io_bresp ;
wire [31:0] _CLINT_io_rdata ;
wire [1:0] _CLINT_io_rresp ;
wire [2:0] _EXU_io_LSUIn_bits_memOp ;
wire [31:0] _EXU_io_LSUIn_bits_raddr ;
wire [31:0] _EXU_io_LSUIn_bits_waddr ;
wire [31:0] _EXU_io_LSUIn_bits_wdata ;
wire [31:0] _EXU_io_out_bits_aluOut ;
wire [1:0] _EXU_io_out_bits_control_wbSrc ;
wire [31:0] _EXU_io_out_bits_csrOut ;
wire [31:0] _EXU_io_out_bits_memOut ;
wire [31:0] _EXU_io_out_bits_pcCom ;
wire [4:0] _EXU_io_out_bits_wa ;
wire [3:0] _IDU_io_RegFileAccess_ra1 ;
wire [3:0] _IDU_io_RegFileAccess_ra2 ;
wire [1:0] _IDU_io_out_bits_control_aluBSrc ;
wire [3:0] _IDU_io_out_bits_control_aluCtr ;
wire [2:0] _IDU_io_out_bits_control_brType ;
wire [2:0] _IDU_io_out_bits_control_csrCtr ;
wire [2:0] _IDU_io_out_bits_control_memOp ;
wire [1:0] _IDU_io_out_bits_control_wbSrc ;
wire [31:0] _IDU_io_out_bits_imm ;
wire [31:0] _IDU_io_out_bits_pc ;
wire [31:0] _IDU_io_out_bits_rd1 ;
wire [31:0] _IDU_io_out_bits_rd2 ;
wire [31:0] _IDU_io_out_bits_uimm ;
wire [4:0] _IDU_io_out_bits_wa ;
wire [31:0] _IFU_io_master_araddr ;
wire [31:0] _IFU_io_out_bits_instruction ;
wire [31:0] _IFU_io_out_bits_pc ;
wire [31:0] _LSU_io_master_araddr ;
wire [2:0] _LSU_io_master_arsize ;
wire [31:0] _LSU_io_master_awaddr ;
wire [2:0] _LSU_io_master_awsize ;
wire [31:0] _LSU_io_master_wdata ;
wire [3:0] _LSU_io_master_wstrb ;
wire [31:0] _LSU_io_out_bits_rdata ;
wire [31:0] _RegFile_io_rd1 ;
wire [31:0] _RegFile_io_rd2 ;
wire [3:0] _WBU_io_RegFileAccess_wa ;
wire [31:0] _WBU_io_RegFileAccess_wd ;
wire [31:0] _WBU_io_out_bits_nextPc ;
wire [31:0] io_master_araddr ;
wire [1:0] io_master_arburst ;
wire [3:0] io_master_arid ;
wire [7:0] io_master_arlen ;
wire [2:0] io_master_arsize ;
wire [31:0] io_master_awaddr ;
wire [1:0] io_master_awburst ;
wire [3:0] io_master_awid ;
wire [7:0] io_master_awlen ;
wire [2:0] io_master_awsize ;
wire [3:0] io_master_bid ;
wire [1:0] io_master_bresp ;
wire [31:0] io_master_rdata ;
wire [3:0] io_master_rid ;
wire [1:0] io_master_rresp ;
wire [31:0] io_master_wdata ;
wire [3:0] io_master_wstrb ;
wire [31:0] io_slave_araddr ;
wire [1:0] io_slave_arburst ;
wire [3:0] io_slave_arid ;
wire [7:0] io_slave_arlen ;
wire [2:0] io_slave_arsize ;
wire [31:0] io_slave_awaddr ;
wire [1:0] io_slave_awburst ;
wire [3:0] io_slave_awid ;
wire [7:0] io_slave_awlen ;
wire [2:0] io_slave_awsize ;
wire [3:0] io_slave_bid ;
wire [1:0] io_slave_bresp ;
wire [31:0] io_slave_rdata ;
wire [3:0] io_slave_rid ;
wire [1:0] io_slave_rresp ;
wire [31:0] io_slave_wdata ;
wire [3:0] io_slave_wstrb ;
wire [1:0] \AXI4Interconnect/state ;
wire [63:0] \CLINT/mtime ;
wire [31:0] \CLINT/readAddr ;
wire [2:0] \CLINT/state ;
wire [31:0] \EXU/casez_tmp_0 ;
wire [1:0] \EXU/in_control_aluBSrc ;
wire [3:0] \EXU/in_control_aluCtr ;
wire [2:0] \EXU/in_control_brType ;
wire [2:0] \EXU/in_control_csrCtr ;
wire [31:0] \EXU/in_imm ;
wire [31:0] \EXU/in_pc ;
wire [31:0] \EXU/in_rd1 ;
wire [31:0] \EXU/in_uimm ;
wire [1:0] \EXU/state ;
wire [31:0] \EXU/ALU/_adder_io_result ;
wire [2:0] \EXU/ALU/_aluControl_io_aluSel ;
wire [31:0] \EXU/ALU/_barrelShift_io_out ;
wire [31:0] \EXU/CSRControl/csrs_0_2 ;
wire [31:0] \EXU/CSRControl/csrs_2_2 ;
wire [31:0] \EXU/CSRControl/csrs_3_2 ;
wire [31:0] \EXU/CSRControl/csrs_4_2 ;
wire [1:0] \EXU/CSRControl/priv ;
wire [2:0] \IDU/_Control_io_immType ;
wire [1:0] \IFU/state ;
wire [2:0] \LSU/in_memOp ;
wire [31:0] \LSU/in_wdata ;
wire [2:0] \LSU/state ;
wire [31:0] \RegFile/reg_0 ;
wire [31:0] \RegFile/reg_10 ;
wire [31:0] \RegFile/reg_11 ;
wire [31:0] \RegFile/reg_12 ;
wire [31:0] \RegFile/reg_13 ;
wire [31:0] \RegFile/reg_14 ;
wire [31:0] \RegFile/reg_15 ;
wire [31:0] \RegFile/reg_1 ;
wire [31:0] \RegFile/reg_2 ;
wire [31:0] \RegFile/reg_3 ;
wire [31:0] \RegFile/reg_4 ;
wire [31:0] \RegFile/reg_5 ;
wire [31:0] \RegFile/reg_6 ;
wire [31:0] \RegFile/reg_7 ;
wire [31:0] \RegFile/reg_8 ;
wire [31:0] \RegFile/reg_9 ;


LOGIC0_X1 _01_ ( .Z(_00_ ) );
BUF_X1 _02_ ( .A(fanout_net_1 ), .Z(\io_master_arid [0] ) );
BUF_X1 _03_ ( .A(fanout_net_1 ), .Z(\io_master_arid [1] ) );
BUF_X1 _04_ ( .A(fanout_net_1 ), .Z(\io_master_arid [2] ) );
BUF_X1 _05_ ( .A(fanout_net_1 ), .Z(\io_master_arid [3] ) );
BUF_X1 _06_ ( .A(fanout_net_1 ), .Z(\io_master_arlen [0] ) );
BUF_X1 _07_ ( .A(fanout_net_1 ), .Z(\io_master_arlen [1] ) );
BUF_X1 _08_ ( .A(fanout_net_1 ), .Z(\io_master_arlen [2] ) );
BUF_X1 _09_ ( .A(fanout_net_1 ), .Z(\io_master_arlen [3] ) );
BUF_X1 _10_ ( .A(fanout_net_1 ), .Z(\io_master_arlen [4] ) );
BUF_X1 _11_ ( .A(fanout_net_1 ), .Z(\io_master_arlen [5] ) );
BUF_X1 _12_ ( .A(fanout_net_1 ), .Z(\io_master_arlen [6] ) );
BUF_X1 _13_ ( .A(fanout_net_1 ), .Z(\io_master_arlen [7] ) );
BUF_X1 _14_ ( .A(fanout_net_1 ), .Z(\io_master_awid [0] ) );
BUF_X1 _15_ ( .A(fanout_net_1 ), .Z(\io_master_awid [1] ) );
BUF_X1 _16_ ( .A(fanout_net_1 ), .Z(\io_master_awid [2] ) );
BUF_X1 _17_ ( .A(fanout_net_1 ), .Z(\io_master_awid [3] ) );
BUF_X1 _18_ ( .A(fanout_net_1 ), .Z(\io_master_awlen [0] ) );
BUF_X1 _19_ ( .A(fanout_net_1 ), .Z(\io_master_awlen [1] ) );
BUF_X1 _20_ ( .A(fanout_net_1 ), .Z(\io_master_awlen [2] ) );
BUF_X1 _21_ ( .A(fanout_net_1 ), .Z(\io_master_awlen [3] ) );
BUF_X1 _22_ ( .A(fanout_net_1 ), .Z(\io_master_awlen [4] ) );
BUF_X1 _23_ ( .A(fanout_net_1 ), .Z(\io_master_awlen [5] ) );
BUF_X1 _24_ ( .A(fanout_net_1 ), .Z(\io_master_awlen [6] ) );
BUF_X1 _25_ ( .A(fanout_net_1 ), .Z(\io_master_awlen [7] ) );
BUF_X1 _26_ ( .A(fanout_net_1 ), .Z(io_slave_arready ) );
BUF_X1 _27_ ( .A(fanout_net_1 ), .Z(io_slave_awready ) );
BUF_X1 _28_ ( .A(fanout_net_1 ), .Z(\io_slave_bid [0] ) );
BUF_X1 _29_ ( .A(fanout_net_1 ), .Z(\io_slave_bid [1] ) );
BUF_X1 _30_ ( .A(fanout_net_1 ), .Z(\io_slave_bid [2] ) );
BUF_X1 _31_ ( .A(fanout_net_1 ), .Z(\io_slave_bid [3] ) );
BUF_X1 _32_ ( .A(fanout_net_2 ), .Z(\io_slave_bresp [0] ) );
BUF_X1 _33_ ( .A(fanout_net_2 ), .Z(\io_slave_bresp [1] ) );
BUF_X1 _34_ ( .A(fanout_net_2 ), .Z(io_slave_bvalid ) );
BUF_X1 _35_ ( .A(fanout_net_2 ), .Z(\io_slave_rdata [0] ) );
BUF_X1 _36_ ( .A(fanout_net_2 ), .Z(\io_slave_rdata [1] ) );
BUF_X1 _37_ ( .A(fanout_net_2 ), .Z(\io_slave_rdata [2] ) );
BUF_X1 _38_ ( .A(fanout_net_2 ), .Z(\io_slave_rdata [3] ) );
BUF_X1 _39_ ( .A(fanout_net_2 ), .Z(\io_slave_rdata [4] ) );
BUF_X1 _40_ ( .A(fanout_net_2 ), .Z(\io_slave_rdata [5] ) );
BUF_X1 _41_ ( .A(fanout_net_2 ), .Z(\io_slave_rdata [6] ) );
BUF_X1 _42_ ( .A(fanout_net_2 ), .Z(\io_slave_rdata [7] ) );
BUF_X1 _43_ ( .A(fanout_net_2 ), .Z(\io_slave_rdata [8] ) );
BUF_X1 _44_ ( .A(fanout_net_2 ), .Z(\io_slave_rdata [9] ) );
BUF_X1 _45_ ( .A(fanout_net_2 ), .Z(\io_slave_rdata [10] ) );
BUF_X1 _46_ ( .A(fanout_net_2 ), .Z(\io_slave_rdata [11] ) );
BUF_X1 _47_ ( .A(fanout_net_2 ), .Z(\io_slave_rdata [12] ) );
BUF_X1 _48_ ( .A(fanout_net_2 ), .Z(\io_slave_rdata [13] ) );
BUF_X1 _49_ ( .A(fanout_net_2 ), .Z(\io_slave_rdata [14] ) );
BUF_X1 _50_ ( .A(fanout_net_2 ), .Z(\io_slave_rdata [15] ) );
BUF_X1 _51_ ( .A(fanout_net_2 ), .Z(\io_slave_rdata [16] ) );
BUF_X1 _52_ ( .A(fanout_net_2 ), .Z(\io_slave_rdata [17] ) );
BUF_X1 _53_ ( .A(fanout_net_2 ), .Z(\io_slave_rdata [18] ) );
BUF_X1 _54_ ( .A(fanout_net_2 ), .Z(\io_slave_rdata [19] ) );
BUF_X1 _55_ ( .A(fanout_net_2 ), .Z(\io_slave_rdata [20] ) );
BUF_X1 _56_ ( .A(fanout_net_2 ), .Z(\io_slave_rdata [21] ) );
BUF_X1 _57_ ( .A(fanout_net_2 ), .Z(\io_slave_rdata [22] ) );
BUF_X1 _58_ ( .A(fanout_net_2 ), .Z(\io_slave_rdata [23] ) );
BUF_X1 _59_ ( .A(fanout_net_2 ), .Z(\io_slave_rdata [24] ) );
BUF_X1 _60_ ( .A(fanout_net_2 ), .Z(\io_slave_rdata [25] ) );
BUF_X1 _61_ ( .A(fanout_net_2 ), .Z(\io_slave_rdata [26] ) );
BUF_X1 _62_ ( .A(_00_ ), .Z(\io_slave_rdata [27] ) );
BUF_X1 _63_ ( .A(_00_ ), .Z(\io_slave_rdata [28] ) );
BUF_X1 _64_ ( .A(_00_ ), .Z(\io_slave_rdata [29] ) );
BUF_X1 _65_ ( .A(_00_ ), .Z(\io_slave_rdata [30] ) );
BUF_X1 _66_ ( .A(_00_ ), .Z(\io_slave_rdata [31] ) );
BUF_X1 _67_ ( .A(_00_ ), .Z(\io_slave_rid [0] ) );
BUF_X1 _68_ ( .A(_00_ ), .Z(\io_slave_rid [1] ) );
BUF_X1 _69_ ( .A(_00_ ), .Z(\io_slave_rid [2] ) );
BUF_X1 _70_ ( .A(_00_ ), .Z(\io_slave_rid [3] ) );
BUF_X1 _71_ ( .A(_00_ ), .Z(io_slave_rlast ) );
BUF_X1 _72_ ( .A(_00_ ), .Z(\io_slave_rresp [0] ) );
BUF_X1 _73_ ( .A(_00_ ), .Z(\io_slave_rresp [1] ) );
BUF_X1 _74_ ( .A(_00_ ), .Z(io_slave_rvalid ) );
BUF_X1 _75_ ( .A(_00_ ), .Z(io_slave_wready ) );
AND2_X1 \AXI4Interconnect/_0881_ ( .A1(\AXI4Interconnect/_0486_ ), .A2(fanout_net_5 ), .ZN(\AXI4Interconnect/_0606_ ) );
INV_X4 \AXI4Interconnect/_0882_ ( .A(fanout_net_5 ), .ZN(\AXI4Interconnect/_0607_ ) );
BUF_X4 \AXI4Interconnect/_0883_ ( .A(\AXI4Interconnect/_0607_ ), .Z(\AXI4Interconnect/_0608_ ) );
AOI21_X1 \AXI4Interconnect/_0884_ ( .A(\AXI4Interconnect/_0606_ ), .B1(\AXI4Interconnect/_0338_ ), .B2(\AXI4Interconnect/_0608_ ), .ZN(\AXI4Interconnect/_0609_ ) );
NOR2_X4 \AXI4Interconnect/_0885_ ( .A1(\AXI4Interconnect/_0873_ ), .A2(\AXI4Interconnect/_0872_ ), .ZN(\AXI4Interconnect/_0610_ ) );
BUF_X8 \AXI4Interconnect/_0886_ ( .A(\AXI4Interconnect/_0610_ ), .Z(\AXI4Interconnect/_0611_ ) );
INV_X1 \AXI4Interconnect/_0887_ ( .A(fanout_net_3 ), .ZN(\AXI4Interconnect/_0612_ ) );
OR2_X1 \AXI4Interconnect/_0888_ ( .A1(\AXI4Interconnect/_0611_ ), .A2(\AXI4Interconnect/_0612_ ), .ZN(\AXI4Interconnect/_0613_ ) );
BUF_X4 \AXI4Interconnect/_0889_ ( .A(\AXI4Interconnect/_0613_ ), .Z(\AXI4Interconnect/_0614_ ) );
BUF_X4 \AXI4Interconnect/_0890_ ( .A(\AXI4Interconnect/_0614_ ), .Z(\AXI4Interconnect/_0615_ ) );
NOR2_X1 \AXI4Interconnect/_0891_ ( .A1(\AXI4Interconnect/_0609_ ), .A2(\AXI4Interconnect/_0615_ ), .ZN(\AXI4Interconnect/_0077_ ) );
AND2_X1 \AXI4Interconnect/_0892_ ( .A1(fanout_net_5 ), .A2(\AXI4Interconnect/_0487_ ), .ZN(\AXI4Interconnect/_0616_ ) );
BUF_X2 \AXI4Interconnect/_0893_ ( .A(\AXI4Interconnect/_0607_ ), .Z(\AXI4Interconnect/_0617_ ) );
BUF_X4 \AXI4Interconnect/_0894_ ( .A(\AXI4Interconnect/_0617_ ), .Z(\AXI4Interconnect/_0618_ ) );
AOI21_X1 \AXI4Interconnect/_0895_ ( .A(\AXI4Interconnect/_0616_ ), .B1(\AXI4Interconnect/_0618_ ), .B2(\AXI4Interconnect/_0339_ ), .ZN(\AXI4Interconnect/_0619_ ) );
NOR2_X1 \AXI4Interconnect/_0896_ ( .A1(\AXI4Interconnect/_0619_ ), .A2(\AXI4Interconnect/_0615_ ), .ZN(\AXI4Interconnect/_0078_ ) );
AND2_X1 \AXI4Interconnect/_0897_ ( .A1(fanout_net_5 ), .A2(\AXI4Interconnect/_0453_ ), .ZN(\AXI4Interconnect/_0620_ ) );
AOI21_X1 \AXI4Interconnect/_0898_ ( .A(\AXI4Interconnect/_0620_ ), .B1(\AXI4Interconnect/_0618_ ), .B2(\AXI4Interconnect/_0305_ ), .ZN(\AXI4Interconnect/_0621_ ) );
NOR2_X1 \AXI4Interconnect/_0899_ ( .A1(\AXI4Interconnect/_0621_ ), .A2(\AXI4Interconnect/_0615_ ), .ZN(\AXI4Interconnect/_0044_ ) );
BUF_X4 \AXI4Interconnect/_0900_ ( .A(\AXI4Interconnect/_0607_ ), .Z(\AXI4Interconnect/_0622_ ) );
OR2_X1 \AXI4Interconnect/_0901_ ( .A1(\AXI4Interconnect/_0622_ ), .A2(\AXI4Interconnect/_0464_ ), .ZN(\AXI4Interconnect/_0623_ ) );
OAI21_X1 \AXI4Interconnect/_0902_ ( .A(\AXI4Interconnect/_0623_ ), .B1(fanout_net_5 ), .B2(\AXI4Interconnect/_0316_ ), .ZN(\AXI4Interconnect/_0624_ ) );
NOR2_X1 \AXI4Interconnect/_0903_ ( .A1(\AXI4Interconnect/_0624_ ), .A2(\AXI4Interconnect/_0615_ ), .ZN(\AXI4Interconnect/_0055_ ) );
OR2_X1 \AXI4Interconnect/_0904_ ( .A1(fanout_net_5 ), .A2(\AXI4Interconnect/_0327_ ), .ZN(\AXI4Interconnect/_0625_ ) );
OAI21_X1 \AXI4Interconnect/_0905_ ( .A(\AXI4Interconnect/_0625_ ), .B1(\AXI4Interconnect/_0608_ ), .B2(\AXI4Interconnect/_0475_ ), .ZN(\AXI4Interconnect/_0626_ ) );
NOR2_X1 \AXI4Interconnect/_0906_ ( .A1(\AXI4Interconnect/_0626_ ), .A2(\AXI4Interconnect/_0615_ ), .ZN(\AXI4Interconnect/_0066_ ) );
AND2_X1 \AXI4Interconnect/_0907_ ( .A1(fanout_net_5 ), .A2(\AXI4Interconnect/_0478_ ), .ZN(\AXI4Interconnect/_0627_ ) );
AOI21_X1 \AXI4Interconnect/_0908_ ( .A(\AXI4Interconnect/_0627_ ), .B1(\AXI4Interconnect/_0618_ ), .B2(\AXI4Interconnect/_0330_ ), .ZN(\AXI4Interconnect/_0628_ ) );
NOR2_X1 \AXI4Interconnect/_0909_ ( .A1(\AXI4Interconnect/_0628_ ), .A2(\AXI4Interconnect/_0615_ ), .ZN(\AXI4Interconnect/_0069_ ) );
OR2_X1 \AXI4Interconnect/_0910_ ( .A1(\AXI4Interconnect/_0622_ ), .A2(\AXI4Interconnect/_0479_ ), .ZN(\AXI4Interconnect/_0629_ ) );
OAI21_X1 \AXI4Interconnect/_0911_ ( .A(\AXI4Interconnect/_0629_ ), .B1(fanout_net_5 ), .B2(\AXI4Interconnect/_0331_ ), .ZN(\AXI4Interconnect/_0630_ ) );
NOR2_X1 \AXI4Interconnect/_0912_ ( .A1(\AXI4Interconnect/_0630_ ), .A2(\AXI4Interconnect/_0615_ ), .ZN(\AXI4Interconnect/_0070_ ) );
AND2_X1 \AXI4Interconnect/_0913_ ( .A1(fanout_net_5 ), .A2(\AXI4Interconnect/_0480_ ), .ZN(\AXI4Interconnect/_0631_ ) );
BUF_X4 \AXI4Interconnect/_0914_ ( .A(\AXI4Interconnect/_0617_ ), .Z(\AXI4Interconnect/_0632_ ) );
AOI21_X1 \AXI4Interconnect/_0915_ ( .A(\AXI4Interconnect/_0631_ ), .B1(\AXI4Interconnect/_0632_ ), .B2(\AXI4Interconnect/_0332_ ), .ZN(\AXI4Interconnect/_0633_ ) );
NOR2_X1 \AXI4Interconnect/_0916_ ( .A1(\AXI4Interconnect/_0633_ ), .A2(\AXI4Interconnect/_0615_ ), .ZN(\AXI4Interconnect/_0071_ ) );
AND2_X1 \AXI4Interconnect/_0917_ ( .A1(fanout_net_5 ), .A2(\AXI4Interconnect/_0481_ ), .ZN(\AXI4Interconnect/_0634_ ) );
AOI21_X1 \AXI4Interconnect/_0918_ ( .A(\AXI4Interconnect/_0634_ ), .B1(\AXI4Interconnect/_0632_ ), .B2(\AXI4Interconnect/_0333_ ), .ZN(\AXI4Interconnect/_0635_ ) );
NOR2_X1 \AXI4Interconnect/_0919_ ( .A1(\AXI4Interconnect/_0635_ ), .A2(\AXI4Interconnect/_0615_ ), .ZN(\AXI4Interconnect/_0072_ ) );
OR2_X1 \AXI4Interconnect/_0920_ ( .A1(\AXI4Interconnect/_0622_ ), .A2(\AXI4Interconnect/_0482_ ), .ZN(\AXI4Interconnect/_0636_ ) );
OAI21_X1 \AXI4Interconnect/_0921_ ( .A(\AXI4Interconnect/_0636_ ), .B1(fanout_net_5 ), .B2(\AXI4Interconnect/_0334_ ), .ZN(\AXI4Interconnect/_0637_ ) );
NOR2_X1 \AXI4Interconnect/_0922_ ( .A1(\AXI4Interconnect/_0637_ ), .A2(\AXI4Interconnect/_0615_ ), .ZN(\AXI4Interconnect/_0073_ ) );
AND2_X1 \AXI4Interconnect/_0923_ ( .A1(fanout_net_5 ), .A2(\AXI4Interconnect/_0483_ ), .ZN(\AXI4Interconnect/_0638_ ) );
AOI21_X1 \AXI4Interconnect/_0924_ ( .A(\AXI4Interconnect/_0638_ ), .B1(\AXI4Interconnect/_0632_ ), .B2(\AXI4Interconnect/_0335_ ), .ZN(\AXI4Interconnect/_0639_ ) );
BUF_X4 \AXI4Interconnect/_0925_ ( .A(\AXI4Interconnect/_0614_ ), .Z(\AXI4Interconnect/_0640_ ) );
NOR2_X1 \AXI4Interconnect/_0926_ ( .A1(\AXI4Interconnect/_0639_ ), .A2(\AXI4Interconnect/_0640_ ), .ZN(\AXI4Interconnect/_0074_ ) );
AND2_X1 \AXI4Interconnect/_0927_ ( .A1(fanout_net_5 ), .A2(\AXI4Interconnect/_0484_ ), .ZN(\AXI4Interconnect/_0641_ ) );
AOI21_X1 \AXI4Interconnect/_0928_ ( .A(\AXI4Interconnect/_0641_ ), .B1(\AXI4Interconnect/_0632_ ), .B2(\AXI4Interconnect/_0336_ ), .ZN(\AXI4Interconnect/_0642_ ) );
NOR2_X1 \AXI4Interconnect/_0929_ ( .A1(\AXI4Interconnect/_0642_ ), .A2(\AXI4Interconnect/_0640_ ), .ZN(\AXI4Interconnect/_0075_ ) );
OR2_X1 \AXI4Interconnect/_0930_ ( .A1(\AXI4Interconnect/_0622_ ), .A2(\AXI4Interconnect/_0454_ ), .ZN(\AXI4Interconnect/_0643_ ) );
OAI21_X1 \AXI4Interconnect/_0931_ ( .A(\AXI4Interconnect/_0643_ ), .B1(fanout_net_5 ), .B2(\AXI4Interconnect/_0306_ ), .ZN(\AXI4Interconnect/_0644_ ) );
NOR2_X1 \AXI4Interconnect/_0932_ ( .A1(\AXI4Interconnect/_0644_ ), .A2(\AXI4Interconnect/_0640_ ), .ZN(\AXI4Interconnect/_0045_ ) );
AND2_X1 \AXI4Interconnect/_0933_ ( .A1(fanout_net_5 ), .A2(\AXI4Interconnect/_0455_ ), .ZN(\AXI4Interconnect/_0645_ ) );
AOI21_X1 \AXI4Interconnect/_0934_ ( .A(\AXI4Interconnect/_0645_ ), .B1(\AXI4Interconnect/_0632_ ), .B2(\AXI4Interconnect/_0307_ ), .ZN(\AXI4Interconnect/_0646_ ) );
NOR2_X1 \AXI4Interconnect/_0935_ ( .A1(\AXI4Interconnect/_0646_ ), .A2(\AXI4Interconnect/_0640_ ), .ZN(\AXI4Interconnect/_0046_ ) );
AND2_X1 \AXI4Interconnect/_0936_ ( .A1(fanout_net_5 ), .A2(\AXI4Interconnect/_0456_ ), .ZN(\AXI4Interconnect/_0647_ ) );
AOI21_X1 \AXI4Interconnect/_0937_ ( .A(\AXI4Interconnect/_0647_ ), .B1(\AXI4Interconnect/_0632_ ), .B2(\AXI4Interconnect/_0308_ ), .ZN(\AXI4Interconnect/_0648_ ) );
NOR2_X1 \AXI4Interconnect/_0938_ ( .A1(\AXI4Interconnect/_0648_ ), .A2(\AXI4Interconnect/_0640_ ), .ZN(\AXI4Interconnect/_0047_ ) );
OR2_X1 \AXI4Interconnect/_0939_ ( .A1(\AXI4Interconnect/_0622_ ), .A2(\AXI4Interconnect/_0457_ ), .ZN(\AXI4Interconnect/_0649_ ) );
OAI21_X1 \AXI4Interconnect/_0940_ ( .A(\AXI4Interconnect/_0649_ ), .B1(fanout_net_5 ), .B2(\AXI4Interconnect/_0309_ ), .ZN(\AXI4Interconnect/_0650_ ) );
NOR2_X1 \AXI4Interconnect/_0941_ ( .A1(\AXI4Interconnect/_0650_ ), .A2(\AXI4Interconnect/_0640_ ), .ZN(\AXI4Interconnect/_0048_ ) );
OR2_X1 \AXI4Interconnect/_0942_ ( .A1(\AXI4Interconnect/_0622_ ), .A2(\AXI4Interconnect/_0458_ ), .ZN(\AXI4Interconnect/_0651_ ) );
OAI21_X1 \AXI4Interconnect/_0943_ ( .A(\AXI4Interconnect/_0651_ ), .B1(fanout_net_5 ), .B2(\AXI4Interconnect/_0310_ ), .ZN(\AXI4Interconnect/_0652_ ) );
NOR2_X1 \AXI4Interconnect/_0944_ ( .A1(\AXI4Interconnect/_0652_ ), .A2(\AXI4Interconnect/_0640_ ), .ZN(\AXI4Interconnect/_0049_ ) );
OR2_X1 \AXI4Interconnect/_0945_ ( .A1(\AXI4Interconnect/_0617_ ), .A2(\AXI4Interconnect/_0459_ ), .ZN(\AXI4Interconnect/_0653_ ) );
OAI21_X1 \AXI4Interconnect/_0946_ ( .A(\AXI4Interconnect/_0653_ ), .B1(fanout_net_5 ), .B2(\AXI4Interconnect/_0311_ ), .ZN(\AXI4Interconnect/_0654_ ) );
NOR2_X1 \AXI4Interconnect/_0947_ ( .A1(\AXI4Interconnect/_0654_ ), .A2(\AXI4Interconnect/_0640_ ), .ZN(\AXI4Interconnect/_0050_ ) );
AND2_X1 \AXI4Interconnect/_0948_ ( .A1(\AXI4Interconnect/_0617_ ), .A2(\AXI4Interconnect/_0312_ ), .ZN(\AXI4Interconnect/_0655_ ) );
AOI21_X1 \AXI4Interconnect/_0949_ ( .A(\AXI4Interconnect/_0655_ ), .B1(fanout_net_5 ), .B2(\AXI4Interconnect/_0460_ ), .ZN(\AXI4Interconnect/_0656_ ) );
NOR2_X1 \AXI4Interconnect/_0950_ ( .A1(\AXI4Interconnect/_0656_ ), .A2(\AXI4Interconnect/_0640_ ), .ZN(\AXI4Interconnect/_0051_ ) );
OR2_X1 \AXI4Interconnect/_0951_ ( .A1(\AXI4Interconnect/_0617_ ), .A2(\AXI4Interconnect/_0461_ ), .ZN(\AXI4Interconnect/_0657_ ) );
OAI21_X1 \AXI4Interconnect/_0952_ ( .A(\AXI4Interconnect/_0657_ ), .B1(fanout_net_5 ), .B2(\AXI4Interconnect/_0313_ ), .ZN(\AXI4Interconnect/_0658_ ) );
NOR2_X1 \AXI4Interconnect/_0953_ ( .A1(\AXI4Interconnect/_0658_ ), .A2(\AXI4Interconnect/_0640_ ), .ZN(\AXI4Interconnect/_0052_ ) );
AND2_X1 \AXI4Interconnect/_0954_ ( .A1(fanout_net_5 ), .A2(\AXI4Interconnect/_0462_ ), .ZN(\AXI4Interconnect/_0659_ ) );
AOI21_X1 \AXI4Interconnect/_0955_ ( .A(\AXI4Interconnect/_0659_ ), .B1(\AXI4Interconnect/_0632_ ), .B2(\AXI4Interconnect/_0314_ ), .ZN(\AXI4Interconnect/_0660_ ) );
BUF_X4 \AXI4Interconnect/_0956_ ( .A(\AXI4Interconnect/_0614_ ), .Z(\AXI4Interconnect/_0661_ ) );
NOR2_X1 \AXI4Interconnect/_0957_ ( .A1(\AXI4Interconnect/_0660_ ), .A2(\AXI4Interconnect/_0661_ ), .ZN(\AXI4Interconnect/_0053_ ) );
OR2_X1 \AXI4Interconnect/_0958_ ( .A1(\AXI4Interconnect/_0617_ ), .A2(\AXI4Interconnect/_0463_ ), .ZN(\AXI4Interconnect/_0662_ ) );
OAI21_X1 \AXI4Interconnect/_0959_ ( .A(\AXI4Interconnect/_0662_ ), .B1(fanout_net_5 ), .B2(\AXI4Interconnect/_0315_ ), .ZN(\AXI4Interconnect/_0663_ ) );
NOR2_X1 \AXI4Interconnect/_0960_ ( .A1(\AXI4Interconnect/_0663_ ), .A2(\AXI4Interconnect/_0661_ ), .ZN(\AXI4Interconnect/_0054_ ) );
AND2_X1 \AXI4Interconnect/_0961_ ( .A1(fanout_net_5 ), .A2(\AXI4Interconnect/_0465_ ), .ZN(\AXI4Interconnect/_0664_ ) );
AOI21_X1 \AXI4Interconnect/_0962_ ( .A(\AXI4Interconnect/_0664_ ), .B1(\AXI4Interconnect/_0632_ ), .B2(\AXI4Interconnect/_0317_ ), .ZN(\AXI4Interconnect/_0665_ ) );
NOR2_X1 \AXI4Interconnect/_0963_ ( .A1(\AXI4Interconnect/_0665_ ), .A2(\AXI4Interconnect/_0661_ ), .ZN(\AXI4Interconnect/_0056_ ) );
AND2_X1 \AXI4Interconnect/_0964_ ( .A1(fanout_net_5 ), .A2(\AXI4Interconnect/_0466_ ), .ZN(\AXI4Interconnect/_0666_ ) );
AOI21_X1 \AXI4Interconnect/_0965_ ( .A(\AXI4Interconnect/_0666_ ), .B1(\AXI4Interconnect/_0632_ ), .B2(\AXI4Interconnect/_0318_ ), .ZN(\AXI4Interconnect/_0667_ ) );
NOR2_X1 \AXI4Interconnect/_0966_ ( .A1(\AXI4Interconnect/_0667_ ), .A2(\AXI4Interconnect/_0661_ ), .ZN(\AXI4Interconnect/_0057_ ) );
AND2_X1 \AXI4Interconnect/_0967_ ( .A1(fanout_net_5 ), .A2(\AXI4Interconnect/_0467_ ), .ZN(\AXI4Interconnect/_0668_ ) );
AOI21_X1 \AXI4Interconnect/_0968_ ( .A(\AXI4Interconnect/_0668_ ), .B1(\AXI4Interconnect/_0632_ ), .B2(\AXI4Interconnect/_0319_ ), .ZN(\AXI4Interconnect/_0669_ ) );
NOR2_X1 \AXI4Interconnect/_0969_ ( .A1(\AXI4Interconnect/_0669_ ), .A2(\AXI4Interconnect/_0661_ ), .ZN(\AXI4Interconnect/_0058_ ) );
AND2_X1 \AXI4Interconnect/_0970_ ( .A1(fanout_net_5 ), .A2(\AXI4Interconnect/_0468_ ), .ZN(\AXI4Interconnect/_0670_ ) );
AOI21_X1 \AXI4Interconnect/_0971_ ( .A(\AXI4Interconnect/_0670_ ), .B1(\AXI4Interconnect/_0608_ ), .B2(\AXI4Interconnect/_0320_ ), .ZN(\AXI4Interconnect/_0671_ ) );
NOR2_X1 \AXI4Interconnect/_0972_ ( .A1(\AXI4Interconnect/_0671_ ), .A2(\AXI4Interconnect/_0661_ ), .ZN(\AXI4Interconnect/_0059_ ) );
AND2_X1 \AXI4Interconnect/_0973_ ( .A1(fanout_net_5 ), .A2(\AXI4Interconnect/_0469_ ), .ZN(\AXI4Interconnect/_0672_ ) );
AOI21_X1 \AXI4Interconnect/_0974_ ( .A(\AXI4Interconnect/_0672_ ), .B1(\AXI4Interconnect/_0608_ ), .B2(\AXI4Interconnect/_0321_ ), .ZN(\AXI4Interconnect/_0673_ ) );
NOR2_X1 \AXI4Interconnect/_0975_ ( .A1(\AXI4Interconnect/_0673_ ), .A2(\AXI4Interconnect/_0661_ ), .ZN(\AXI4Interconnect/_0060_ ) );
AND2_X1 \AXI4Interconnect/_0976_ ( .A1(fanout_net_5 ), .A2(\AXI4Interconnect/_0470_ ), .ZN(\AXI4Interconnect/_0674_ ) );
AOI21_X1 \AXI4Interconnect/_0977_ ( .A(\AXI4Interconnect/_0674_ ), .B1(\AXI4Interconnect/_0608_ ), .B2(\AXI4Interconnect/_0322_ ), .ZN(\AXI4Interconnect/_0675_ ) );
NOR2_X1 \AXI4Interconnect/_0978_ ( .A1(\AXI4Interconnect/_0675_ ), .A2(\AXI4Interconnect/_0661_ ), .ZN(\AXI4Interconnect/_0061_ ) );
OR2_X1 \AXI4Interconnect/_0979_ ( .A1(\AXI4Interconnect/_0617_ ), .A2(\AXI4Interconnect/_0471_ ), .ZN(\AXI4Interconnect/_0676_ ) );
OAI21_X1 \AXI4Interconnect/_0980_ ( .A(\AXI4Interconnect/_0676_ ), .B1(fanout_net_5 ), .B2(\AXI4Interconnect/_0323_ ), .ZN(\AXI4Interconnect/_0677_ ) );
NOR2_X1 \AXI4Interconnect/_0981_ ( .A1(\AXI4Interconnect/_0677_ ), .A2(\AXI4Interconnect/_0661_ ), .ZN(\AXI4Interconnect/_0062_ ) );
OR2_X1 \AXI4Interconnect/_0982_ ( .A1(\AXI4Interconnect/_0617_ ), .A2(\AXI4Interconnect/_0472_ ), .ZN(\AXI4Interconnect/_0678_ ) );
OAI21_X1 \AXI4Interconnect/_0983_ ( .A(\AXI4Interconnect/_0678_ ), .B1(\AXI4Interconnect/_0869_ ), .B2(\AXI4Interconnect/_0324_ ), .ZN(\AXI4Interconnect/_0679_ ) );
NOR2_X1 \AXI4Interconnect/_0984_ ( .A1(\AXI4Interconnect/_0679_ ), .A2(\AXI4Interconnect/_0661_ ), .ZN(\AXI4Interconnect/_0063_ ) );
AND2_X1 \AXI4Interconnect/_0985_ ( .A1(\AXI4Interconnect/_0869_ ), .A2(\AXI4Interconnect/_0473_ ), .ZN(\AXI4Interconnect/_0680_ ) );
AOI21_X1 \AXI4Interconnect/_0986_ ( .A(\AXI4Interconnect/_0680_ ), .B1(\AXI4Interconnect/_0608_ ), .B2(\AXI4Interconnect/_0325_ ), .ZN(\AXI4Interconnect/_0681_ ) );
NOR2_X1 \AXI4Interconnect/_0987_ ( .A1(\AXI4Interconnect/_0681_ ), .A2(\AXI4Interconnect/_0614_ ), .ZN(\AXI4Interconnect/_0064_ ) );
OR2_X1 \AXI4Interconnect/_0988_ ( .A1(\AXI4Interconnect/_0617_ ), .A2(\AXI4Interconnect/_0474_ ), .ZN(\AXI4Interconnect/_0682_ ) );
OAI21_X1 \AXI4Interconnect/_0989_ ( .A(\AXI4Interconnect/_0682_ ), .B1(\AXI4Interconnect/_0869_ ), .B2(\AXI4Interconnect/_0326_ ), .ZN(\AXI4Interconnect/_0683_ ) );
NOR2_X1 \AXI4Interconnect/_0990_ ( .A1(\AXI4Interconnect/_0683_ ), .A2(\AXI4Interconnect/_0614_ ), .ZN(\AXI4Interconnect/_0065_ ) );
AND2_X1 \AXI4Interconnect/_0991_ ( .A1(\AXI4Interconnect/_0869_ ), .A2(\AXI4Interconnect/_0476_ ), .ZN(\AXI4Interconnect/_0684_ ) );
AOI21_X1 \AXI4Interconnect/_0992_ ( .A(\AXI4Interconnect/_0684_ ), .B1(\AXI4Interconnect/_0608_ ), .B2(\AXI4Interconnect/_0328_ ), .ZN(\AXI4Interconnect/_0685_ ) );
NOR2_X1 \AXI4Interconnect/_0993_ ( .A1(\AXI4Interconnect/_0685_ ), .A2(\AXI4Interconnect/_0614_ ), .ZN(\AXI4Interconnect/_0067_ ) );
AND2_X1 \AXI4Interconnect/_0994_ ( .A1(\AXI4Interconnect/_0869_ ), .A2(\AXI4Interconnect/_0477_ ), .ZN(\AXI4Interconnect/_0686_ ) );
AOI21_X1 \AXI4Interconnect/_0995_ ( .A(\AXI4Interconnect/_0686_ ), .B1(\AXI4Interconnect/_0608_ ), .B2(\AXI4Interconnect/_0329_ ), .ZN(\AXI4Interconnect/_0687_ ) );
NOR2_X1 \AXI4Interconnect/_0996_ ( .A1(\AXI4Interconnect/_0687_ ), .A2(\AXI4Interconnect/_0614_ ), .ZN(\AXI4Interconnect/_0068_ ) );
MUX2_X1 \AXI4Interconnect/_0997_ ( .A(\AXI4Interconnect/_0302_ ), .B(\AXI4Interconnect/_0450_ ), .S(\AXI4Interconnect/_0869_ ), .Z(\AXI4Interconnect/_0688_ ) );
INV_X32 \AXI4Interconnect/_0998_ ( .A(fanout_net_6 ), .ZN(\AXI4Interconnect/_0689_ ) );
NOR2_X4 \AXI4Interconnect/_0999_ ( .A1(\AXI4Interconnect/_0611_ ), .A2(\AXI4Interconnect/_0689_ ), .ZN(\AXI4Interconnect/_0690_ ) );
AND2_X1 \AXI4Interconnect/_1000_ ( .A1(\AXI4Interconnect/_0688_ ), .A2(\AXI4Interconnect/_0690_ ), .ZN(\AXI4Interconnect/_0155_ ) );
MUX2_X1 \AXI4Interconnect/_1001_ ( .A(\AXI4Interconnect/_0303_ ), .B(\AXI4Interconnect/_0451_ ), .S(\AXI4Interconnect/_0869_ ), .Z(\AXI4Interconnect/_0691_ ) );
AND2_X1 \AXI4Interconnect/_1002_ ( .A1(\AXI4Interconnect/_0691_ ), .A2(\AXI4Interconnect/_0690_ ), .ZN(\AXI4Interconnect/_0156_ ) );
INV_X2 \AXI4Interconnect/_1003_ ( .A(\AXI4Interconnect/_0690_ ), .ZN(\AXI4Interconnect/_0692_ ) );
BUF_X4 \AXI4Interconnect/_1004_ ( .A(\AXI4Interconnect/_0692_ ), .Z(\AXI4Interconnect/_0693_ ) );
NOR2_X1 \AXI4Interconnect/_1005_ ( .A1(\AXI4Interconnect/_0693_ ), .A2(\AXI4Interconnect/_0609_ ), .ZN(\AXI4Interconnect/_0191_ ) );
NOR2_X1 \AXI4Interconnect/_1006_ ( .A1(\AXI4Interconnect/_0693_ ), .A2(\AXI4Interconnect/_0619_ ), .ZN(\AXI4Interconnect/_0192_ ) );
NOR2_X1 \AXI4Interconnect/_1007_ ( .A1(\AXI4Interconnect/_0693_ ), .A2(\AXI4Interconnect/_0621_ ), .ZN(\AXI4Interconnect/_0158_ ) );
BUF_X4 \AXI4Interconnect/_1008_ ( .A(\AXI4Interconnect/_0692_ ), .Z(\AXI4Interconnect/_0694_ ) );
NOR2_X1 \AXI4Interconnect/_1009_ ( .A1(\AXI4Interconnect/_0624_ ), .A2(\AXI4Interconnect/_0694_ ), .ZN(\AXI4Interconnect/_0169_ ) );
NOR2_X1 \AXI4Interconnect/_1010_ ( .A1(\AXI4Interconnect/_0693_ ), .A2(\AXI4Interconnect/_0626_ ), .ZN(\AXI4Interconnect/_0180_ ) );
NOR2_X1 \AXI4Interconnect/_1011_ ( .A1(\AXI4Interconnect/_0693_ ), .A2(\AXI4Interconnect/_0628_ ), .ZN(\AXI4Interconnect/_0183_ ) );
NOR2_X1 \AXI4Interconnect/_1012_ ( .A1(\AXI4Interconnect/_0630_ ), .A2(\AXI4Interconnect/_0694_ ), .ZN(\AXI4Interconnect/_0184_ ) );
NOR2_X1 \AXI4Interconnect/_1013_ ( .A1(\AXI4Interconnect/_0693_ ), .A2(\AXI4Interconnect/_0633_ ), .ZN(\AXI4Interconnect/_0185_ ) );
NOR2_X1 \AXI4Interconnect/_1014_ ( .A1(\AXI4Interconnect/_0693_ ), .A2(\AXI4Interconnect/_0635_ ), .ZN(\AXI4Interconnect/_0186_ ) );
NOR2_X1 \AXI4Interconnect/_1015_ ( .A1(\AXI4Interconnect/_0637_ ), .A2(\AXI4Interconnect/_0694_ ), .ZN(\AXI4Interconnect/_0187_ ) );
NOR2_X1 \AXI4Interconnect/_1016_ ( .A1(\AXI4Interconnect/_0693_ ), .A2(\AXI4Interconnect/_0639_ ), .ZN(\AXI4Interconnect/_0188_ ) );
NOR2_X1 \AXI4Interconnect/_1017_ ( .A1(\AXI4Interconnect/_0693_ ), .A2(\AXI4Interconnect/_0642_ ), .ZN(\AXI4Interconnect/_0189_ ) );
NOR2_X1 \AXI4Interconnect/_1018_ ( .A1(\AXI4Interconnect/_0644_ ), .A2(\AXI4Interconnect/_0694_ ), .ZN(\AXI4Interconnect/_0159_ ) );
NOR2_X1 \AXI4Interconnect/_1019_ ( .A1(\AXI4Interconnect/_0693_ ), .A2(\AXI4Interconnect/_0646_ ), .ZN(\AXI4Interconnect/_0160_ ) );
BUF_X4 \AXI4Interconnect/_1020_ ( .A(\AXI4Interconnect/_0692_ ), .Z(\AXI4Interconnect/_0695_ ) );
NOR2_X1 \AXI4Interconnect/_1021_ ( .A1(\AXI4Interconnect/_0695_ ), .A2(\AXI4Interconnect/_0648_ ), .ZN(\AXI4Interconnect/_0161_ ) );
NOR2_X1 \AXI4Interconnect/_1022_ ( .A1(\AXI4Interconnect/_0650_ ), .A2(\AXI4Interconnect/_0694_ ), .ZN(\AXI4Interconnect/_0162_ ) );
NOR2_X1 \AXI4Interconnect/_1023_ ( .A1(\AXI4Interconnect/_0652_ ), .A2(\AXI4Interconnect/_0694_ ), .ZN(\AXI4Interconnect/_0163_ ) );
NOR2_X1 \AXI4Interconnect/_1024_ ( .A1(\AXI4Interconnect/_0654_ ), .A2(\AXI4Interconnect/_0694_ ), .ZN(\AXI4Interconnect/_0164_ ) );
NOR2_X1 \AXI4Interconnect/_1025_ ( .A1(\AXI4Interconnect/_0656_ ), .A2(\AXI4Interconnect/_0694_ ), .ZN(\AXI4Interconnect/_0165_ ) );
NOR2_X1 \AXI4Interconnect/_1026_ ( .A1(\AXI4Interconnect/_0658_ ), .A2(\AXI4Interconnect/_0694_ ), .ZN(\AXI4Interconnect/_0166_ ) );
NOR2_X1 \AXI4Interconnect/_1027_ ( .A1(\AXI4Interconnect/_0695_ ), .A2(\AXI4Interconnect/_0660_ ), .ZN(\AXI4Interconnect/_0167_ ) );
NOR2_X1 \AXI4Interconnect/_1028_ ( .A1(\AXI4Interconnect/_0663_ ), .A2(\AXI4Interconnect/_0692_ ), .ZN(\AXI4Interconnect/_0168_ ) );
NOR2_X1 \AXI4Interconnect/_1029_ ( .A1(\AXI4Interconnect/_0695_ ), .A2(\AXI4Interconnect/_0665_ ), .ZN(\AXI4Interconnect/_0170_ ) );
NOR2_X1 \AXI4Interconnect/_1030_ ( .A1(\AXI4Interconnect/_0695_ ), .A2(\AXI4Interconnect/_0667_ ), .ZN(\AXI4Interconnect/_0171_ ) );
NOR2_X1 \AXI4Interconnect/_1031_ ( .A1(\AXI4Interconnect/_0695_ ), .A2(\AXI4Interconnect/_0669_ ), .ZN(\AXI4Interconnect/_0172_ ) );
NOR2_X1 \AXI4Interconnect/_1032_ ( .A1(\AXI4Interconnect/_0695_ ), .A2(\AXI4Interconnect/_0671_ ), .ZN(\AXI4Interconnect/_0173_ ) );
NOR2_X1 \AXI4Interconnect/_1033_ ( .A1(\AXI4Interconnect/_0695_ ), .A2(\AXI4Interconnect/_0673_ ), .ZN(\AXI4Interconnect/_0174_ ) );
NOR2_X1 \AXI4Interconnect/_1034_ ( .A1(\AXI4Interconnect/_0695_ ), .A2(\AXI4Interconnect/_0675_ ), .ZN(\AXI4Interconnect/_0175_ ) );
NOR2_X1 \AXI4Interconnect/_1035_ ( .A1(\AXI4Interconnect/_0677_ ), .A2(\AXI4Interconnect/_0692_ ), .ZN(\AXI4Interconnect/_0176_ ) );
NOR2_X1 \AXI4Interconnect/_1036_ ( .A1(\AXI4Interconnect/_0679_ ), .A2(\AXI4Interconnect/_0692_ ), .ZN(\AXI4Interconnect/_0177_ ) );
NOR2_X1 \AXI4Interconnect/_1037_ ( .A1(\AXI4Interconnect/_0695_ ), .A2(\AXI4Interconnect/_0681_ ), .ZN(\AXI4Interconnect/_0178_ ) );
NOR2_X1 \AXI4Interconnect/_1038_ ( .A1(\AXI4Interconnect/_0683_ ), .A2(\AXI4Interconnect/_0692_ ), .ZN(\AXI4Interconnect/_0179_ ) );
NOR2_X1 \AXI4Interconnect/_1039_ ( .A1(\AXI4Interconnect/_0695_ ), .A2(\AXI4Interconnect/_0685_ ), .ZN(\AXI4Interconnect/_0181_ ) );
NOR2_X1 \AXI4Interconnect/_1040_ ( .A1(\AXI4Interconnect/_0694_ ), .A2(\AXI4Interconnect/_0687_ ), .ZN(\AXI4Interconnect/_0182_ ) );
BUF_X4 \AXI4Interconnect/_1041_ ( .A(\AXI4Interconnect/_0611_ ), .Z(\AXI4Interconnect/_0696_ ) );
BUF_X4 \AXI4Interconnect/_1042_ ( .A(\AXI4Interconnect/_0696_ ), .Z(\AXI4Interconnect/_0697_ ) );
BUF_X4 \AXI4Interconnect/_1043_ ( .A(\AXI4Interconnect/_0689_ ), .Z(\AXI4Interconnect/_0698_ ) );
BUF_X4 \AXI4Interconnect/_1044_ ( .A(\AXI4Interconnect/_0698_ ), .Z(\AXI4Interconnect/_0699_ ) );
BUF_X4 \AXI4Interconnect/_1045_ ( .A(\AXI4Interconnect/_0699_ ), .Z(\AXI4Interconnect/_0700_ ) );
INV_X1 \AXI4Interconnect/_1046_ ( .A(\AXI4Interconnect/_0005_ ), .ZN(\AXI4Interconnect/_0701_ ) );
BUF_X4 \AXI4Interconnect/_1047_ ( .A(\AXI4Interconnect/_0701_ ), .Z(\AXI4Interconnect/_0702_ ) );
BUF_X4 \AXI4Interconnect/_1048_ ( .A(\AXI4Interconnect/_0702_ ), .Z(\AXI4Interconnect/_0703_ ) );
INV_X1 \AXI4Interconnect/_1049_ ( .A(\AXI4Interconnect/_0117_ ), .ZN(\AXI4Interconnect/_0704_ ) );
NOR4_X1 \AXI4Interconnect/_1050_ ( .A1(\AXI4Interconnect/_0697_ ), .A2(\AXI4Interconnect/_0700_ ), .A3(\AXI4Interconnect/_0703_ ), .A4(\AXI4Interconnect/_0704_ ), .ZN(\AXI4Interconnect/_0267_ ) );
INV_X1 \AXI4Interconnect/_1051_ ( .A(\AXI4Interconnect/_0128_ ), .ZN(\AXI4Interconnect/_0705_ ) );
NOR4_X1 \AXI4Interconnect/_1052_ ( .A1(\AXI4Interconnect/_0697_ ), .A2(\AXI4Interconnect/_0700_ ), .A3(\AXI4Interconnect/_0703_ ), .A4(\AXI4Interconnect/_0705_ ), .ZN(\AXI4Interconnect/_0278_ ) );
INV_X1 \AXI4Interconnect/_1053_ ( .A(\AXI4Interconnect/_0139_ ), .ZN(\AXI4Interconnect/_0706_ ) );
NOR4_X1 \AXI4Interconnect/_1054_ ( .A1(\AXI4Interconnect/_0697_ ), .A2(\AXI4Interconnect/_0700_ ), .A3(\AXI4Interconnect/_0703_ ), .A4(\AXI4Interconnect/_0706_ ), .ZN(\AXI4Interconnect/_0289_ ) );
INV_X1 \AXI4Interconnect/_1055_ ( .A(\AXI4Interconnect/_0142_ ), .ZN(\AXI4Interconnect/_0707_ ) );
NOR4_X1 \AXI4Interconnect/_1056_ ( .A1(\AXI4Interconnect/_0697_ ), .A2(\AXI4Interconnect/_0700_ ), .A3(\AXI4Interconnect/_0703_ ), .A4(\AXI4Interconnect/_0707_ ), .ZN(\AXI4Interconnect/_0292_ ) );
INV_X1 \AXI4Interconnect/_1057_ ( .A(\AXI4Interconnect/_0143_ ), .ZN(\AXI4Interconnect/_0708_ ) );
NOR4_X1 \AXI4Interconnect/_1058_ ( .A1(\AXI4Interconnect/_0697_ ), .A2(\AXI4Interconnect/_0700_ ), .A3(\AXI4Interconnect/_0703_ ), .A4(\AXI4Interconnect/_0708_ ), .ZN(\AXI4Interconnect/_0293_ ) );
INV_X1 \AXI4Interconnect/_1059_ ( .A(\AXI4Interconnect/_0144_ ), .ZN(\AXI4Interconnect/_0709_ ) );
NOR4_X1 \AXI4Interconnect/_1060_ ( .A1(\AXI4Interconnect/_0697_ ), .A2(\AXI4Interconnect/_0700_ ), .A3(\AXI4Interconnect/_0703_ ), .A4(\AXI4Interconnect/_0709_ ), .ZN(\AXI4Interconnect/_0294_ ) );
INV_X1 \AXI4Interconnect/_1061_ ( .A(\AXI4Interconnect/_0145_ ), .ZN(\AXI4Interconnect/_0710_ ) );
NOR4_X1 \AXI4Interconnect/_1062_ ( .A1(\AXI4Interconnect/_0697_ ), .A2(\AXI4Interconnect/_0700_ ), .A3(\AXI4Interconnect/_0703_ ), .A4(\AXI4Interconnect/_0710_ ), .ZN(\AXI4Interconnect/_0295_ ) );
INV_X1 \AXI4Interconnect/_1063_ ( .A(\AXI4Interconnect/_0146_ ), .ZN(\AXI4Interconnect/_0711_ ) );
NOR4_X1 \AXI4Interconnect/_1064_ ( .A1(\AXI4Interconnect/_0697_ ), .A2(\AXI4Interconnect/_0700_ ), .A3(\AXI4Interconnect/_0703_ ), .A4(\AXI4Interconnect/_0711_ ), .ZN(\AXI4Interconnect/_0296_ ) );
BUF_X4 \AXI4Interconnect/_1065_ ( .A(\AXI4Interconnect/_0698_ ), .Z(\AXI4Interconnect/_0712_ ) );
BUF_X4 \AXI4Interconnect/_1066_ ( .A(\AXI4Interconnect/_0712_ ), .Z(\AXI4Interconnect/_0713_ ) );
INV_X1 \AXI4Interconnect/_1067_ ( .A(\AXI4Interconnect/_0147_ ), .ZN(\AXI4Interconnect/_0714_ ) );
NOR4_X1 \AXI4Interconnect/_1068_ ( .A1(\AXI4Interconnect/_0697_ ), .A2(\AXI4Interconnect/_0713_ ), .A3(\AXI4Interconnect/_0703_ ), .A4(\AXI4Interconnect/_0714_ ), .ZN(\AXI4Interconnect/_0297_ ) );
INV_X1 \AXI4Interconnect/_1069_ ( .A(\AXI4Interconnect/_0148_ ), .ZN(\AXI4Interconnect/_0715_ ) );
NOR4_X1 \AXI4Interconnect/_1070_ ( .A1(\AXI4Interconnect/_0697_ ), .A2(\AXI4Interconnect/_0713_ ), .A3(\AXI4Interconnect/_0703_ ), .A4(\AXI4Interconnect/_0715_ ), .ZN(\AXI4Interconnect/_0298_ ) );
BUF_X4 \AXI4Interconnect/_1071_ ( .A(\AXI4Interconnect/_0696_ ), .Z(\AXI4Interconnect/_0716_ ) );
BUF_X4 \AXI4Interconnect/_1072_ ( .A(\AXI4Interconnect/_0702_ ), .Z(\AXI4Interconnect/_0717_ ) );
INV_X1 \AXI4Interconnect/_1073_ ( .A(\AXI4Interconnect/_0118_ ), .ZN(\AXI4Interconnect/_0718_ ) );
NOR4_X1 \AXI4Interconnect/_1074_ ( .A1(\AXI4Interconnect/_0716_ ), .A2(\AXI4Interconnect/_0713_ ), .A3(\AXI4Interconnect/_0717_ ), .A4(\AXI4Interconnect/_0718_ ), .ZN(\AXI4Interconnect/_0268_ ) );
INV_X1 \AXI4Interconnect/_1075_ ( .A(\AXI4Interconnect/_0119_ ), .ZN(\AXI4Interconnect/_0719_ ) );
NOR4_X1 \AXI4Interconnect/_1076_ ( .A1(\AXI4Interconnect/_0716_ ), .A2(\AXI4Interconnect/_0713_ ), .A3(\AXI4Interconnect/_0717_ ), .A4(\AXI4Interconnect/_0719_ ), .ZN(\AXI4Interconnect/_0269_ ) );
INV_X1 \AXI4Interconnect/_1077_ ( .A(\AXI4Interconnect/_0120_ ), .ZN(\AXI4Interconnect/_0720_ ) );
NOR4_X1 \AXI4Interconnect/_1078_ ( .A1(\AXI4Interconnect/_0716_ ), .A2(\AXI4Interconnect/_0713_ ), .A3(\AXI4Interconnect/_0717_ ), .A4(\AXI4Interconnect/_0720_ ), .ZN(\AXI4Interconnect/_0270_ ) );
INV_X1 \AXI4Interconnect/_1079_ ( .A(\AXI4Interconnect/_0121_ ), .ZN(\AXI4Interconnect/_0721_ ) );
NOR4_X1 \AXI4Interconnect/_1080_ ( .A1(\AXI4Interconnect/_0716_ ), .A2(\AXI4Interconnect/_0713_ ), .A3(\AXI4Interconnect/_0717_ ), .A4(\AXI4Interconnect/_0721_ ), .ZN(\AXI4Interconnect/_0271_ ) );
INV_X1 \AXI4Interconnect/_1081_ ( .A(\AXI4Interconnect/_0122_ ), .ZN(\AXI4Interconnect/_0722_ ) );
NOR4_X1 \AXI4Interconnect/_1082_ ( .A1(\AXI4Interconnect/_0716_ ), .A2(\AXI4Interconnect/_0713_ ), .A3(\AXI4Interconnect/_0717_ ), .A4(\AXI4Interconnect/_0722_ ), .ZN(\AXI4Interconnect/_0272_ ) );
INV_X1 \AXI4Interconnect/_1083_ ( .A(\AXI4Interconnect/_0123_ ), .ZN(\AXI4Interconnect/_0723_ ) );
NOR4_X1 \AXI4Interconnect/_1084_ ( .A1(\AXI4Interconnect/_0716_ ), .A2(\AXI4Interconnect/_0713_ ), .A3(\AXI4Interconnect/_0717_ ), .A4(\AXI4Interconnect/_0723_ ), .ZN(\AXI4Interconnect/_0273_ ) );
INV_X1 \AXI4Interconnect/_1085_ ( .A(\AXI4Interconnect/_0124_ ), .ZN(\AXI4Interconnect/_0724_ ) );
NOR4_X1 \AXI4Interconnect/_1086_ ( .A1(\AXI4Interconnect/_0716_ ), .A2(\AXI4Interconnect/_0713_ ), .A3(\AXI4Interconnect/_0717_ ), .A4(\AXI4Interconnect/_0724_ ), .ZN(\AXI4Interconnect/_0274_ ) );
INV_X1 \AXI4Interconnect/_1087_ ( .A(\AXI4Interconnect/_0125_ ), .ZN(\AXI4Interconnect/_0725_ ) );
NOR4_X1 \AXI4Interconnect/_1088_ ( .A1(\AXI4Interconnect/_0716_ ), .A2(\AXI4Interconnect/_0713_ ), .A3(\AXI4Interconnect/_0717_ ), .A4(\AXI4Interconnect/_0725_ ), .ZN(\AXI4Interconnect/_0275_ ) );
BUF_X4 \AXI4Interconnect/_1089_ ( .A(\AXI4Interconnect/_0712_ ), .Z(\AXI4Interconnect/_0726_ ) );
INV_X1 \AXI4Interconnect/_1090_ ( .A(\AXI4Interconnect/_0126_ ), .ZN(\AXI4Interconnect/_0727_ ) );
NOR4_X1 \AXI4Interconnect/_1091_ ( .A1(\AXI4Interconnect/_0716_ ), .A2(\AXI4Interconnect/_0726_ ), .A3(\AXI4Interconnect/_0717_ ), .A4(\AXI4Interconnect/_0727_ ), .ZN(\AXI4Interconnect/_0276_ ) );
INV_X1 \AXI4Interconnect/_1092_ ( .A(\AXI4Interconnect/_0127_ ), .ZN(\AXI4Interconnect/_0728_ ) );
NOR4_X1 \AXI4Interconnect/_1093_ ( .A1(\AXI4Interconnect/_0716_ ), .A2(\AXI4Interconnect/_0726_ ), .A3(\AXI4Interconnect/_0717_ ), .A4(\AXI4Interconnect/_0728_ ), .ZN(\AXI4Interconnect/_0277_ ) );
BUF_X4 \AXI4Interconnect/_1094_ ( .A(\AXI4Interconnect/_0696_ ), .Z(\AXI4Interconnect/_0729_ ) );
BUF_X4 \AXI4Interconnect/_1095_ ( .A(\AXI4Interconnect/_0702_ ), .Z(\AXI4Interconnect/_0730_ ) );
INV_X1 \AXI4Interconnect/_1096_ ( .A(\AXI4Interconnect/_0129_ ), .ZN(\AXI4Interconnect/_0731_ ) );
NOR4_X1 \AXI4Interconnect/_1097_ ( .A1(\AXI4Interconnect/_0729_ ), .A2(\AXI4Interconnect/_0726_ ), .A3(\AXI4Interconnect/_0730_ ), .A4(\AXI4Interconnect/_0731_ ), .ZN(\AXI4Interconnect/_0279_ ) );
INV_X1 \AXI4Interconnect/_1098_ ( .A(\AXI4Interconnect/_0130_ ), .ZN(\AXI4Interconnect/_0732_ ) );
NOR4_X1 \AXI4Interconnect/_1099_ ( .A1(\AXI4Interconnect/_0729_ ), .A2(\AXI4Interconnect/_0726_ ), .A3(\AXI4Interconnect/_0730_ ), .A4(\AXI4Interconnect/_0732_ ), .ZN(\AXI4Interconnect/_0280_ ) );
INV_X1 \AXI4Interconnect/_1100_ ( .A(\AXI4Interconnect/_0131_ ), .ZN(\AXI4Interconnect/_0733_ ) );
NOR4_X1 \AXI4Interconnect/_1101_ ( .A1(\AXI4Interconnect/_0729_ ), .A2(\AXI4Interconnect/_0726_ ), .A3(\AXI4Interconnect/_0730_ ), .A4(\AXI4Interconnect/_0733_ ), .ZN(\AXI4Interconnect/_0281_ ) );
INV_X1 \AXI4Interconnect/_1102_ ( .A(\AXI4Interconnect/_0132_ ), .ZN(\AXI4Interconnect/_0734_ ) );
NOR4_X1 \AXI4Interconnect/_1103_ ( .A1(\AXI4Interconnect/_0729_ ), .A2(\AXI4Interconnect/_0726_ ), .A3(\AXI4Interconnect/_0730_ ), .A4(\AXI4Interconnect/_0734_ ), .ZN(\AXI4Interconnect/_0282_ ) );
INV_X1 \AXI4Interconnect/_1104_ ( .A(\AXI4Interconnect/_0133_ ), .ZN(\AXI4Interconnect/_0735_ ) );
NOR4_X1 \AXI4Interconnect/_1105_ ( .A1(\AXI4Interconnect/_0729_ ), .A2(\AXI4Interconnect/_0726_ ), .A3(\AXI4Interconnect/_0730_ ), .A4(\AXI4Interconnect/_0735_ ), .ZN(\AXI4Interconnect/_0283_ ) );
INV_X1 \AXI4Interconnect/_1106_ ( .A(\AXI4Interconnect/_0134_ ), .ZN(\AXI4Interconnect/_0736_ ) );
NOR4_X1 \AXI4Interconnect/_1107_ ( .A1(\AXI4Interconnect/_0729_ ), .A2(\AXI4Interconnect/_0726_ ), .A3(\AXI4Interconnect/_0730_ ), .A4(\AXI4Interconnect/_0736_ ), .ZN(\AXI4Interconnect/_0284_ ) );
INV_X1 \AXI4Interconnect/_1108_ ( .A(\AXI4Interconnect/_0135_ ), .ZN(\AXI4Interconnect/_0737_ ) );
NOR4_X1 \AXI4Interconnect/_1109_ ( .A1(\AXI4Interconnect/_0729_ ), .A2(\AXI4Interconnect/_0726_ ), .A3(\AXI4Interconnect/_0730_ ), .A4(\AXI4Interconnect/_0737_ ), .ZN(\AXI4Interconnect/_0285_ ) );
INV_X1 \AXI4Interconnect/_1110_ ( .A(\AXI4Interconnect/_0136_ ), .ZN(\AXI4Interconnect/_0738_ ) );
NOR4_X1 \AXI4Interconnect/_1111_ ( .A1(\AXI4Interconnect/_0729_ ), .A2(\AXI4Interconnect/_0726_ ), .A3(\AXI4Interconnect/_0730_ ), .A4(\AXI4Interconnect/_0738_ ), .ZN(\AXI4Interconnect/_0286_ ) );
BUF_X4 \AXI4Interconnect/_1112_ ( .A(\AXI4Interconnect/_0712_ ), .Z(\AXI4Interconnect/_0739_ ) );
INV_X1 \AXI4Interconnect/_1113_ ( .A(\AXI4Interconnect/_0137_ ), .ZN(\AXI4Interconnect/_0740_ ) );
NOR4_X1 \AXI4Interconnect/_1114_ ( .A1(\AXI4Interconnect/_0729_ ), .A2(\AXI4Interconnect/_0739_ ), .A3(\AXI4Interconnect/_0730_ ), .A4(\AXI4Interconnect/_0740_ ), .ZN(\AXI4Interconnect/_0287_ ) );
INV_X1 \AXI4Interconnect/_1115_ ( .A(\AXI4Interconnect/_0138_ ), .ZN(\AXI4Interconnect/_0741_ ) );
NOR4_X1 \AXI4Interconnect/_1116_ ( .A1(\AXI4Interconnect/_0729_ ), .A2(\AXI4Interconnect/_0739_ ), .A3(\AXI4Interconnect/_0730_ ), .A4(\AXI4Interconnect/_0741_ ), .ZN(\AXI4Interconnect/_0288_ ) );
BUF_X8 \AXI4Interconnect/_1117_ ( .A(\AXI4Interconnect/_0611_ ), .Z(\AXI4Interconnect/_0742_ ) );
BUF_X4 \AXI4Interconnect/_1118_ ( .A(\AXI4Interconnect/_0742_ ), .Z(\AXI4Interconnect/_0743_ ) );
BUF_X4 \AXI4Interconnect/_1119_ ( .A(\AXI4Interconnect/_0702_ ), .Z(\AXI4Interconnect/_0744_ ) );
INV_X1 \AXI4Interconnect/_1120_ ( .A(\AXI4Interconnect/_0140_ ), .ZN(\AXI4Interconnect/_0745_ ) );
NOR4_X1 \AXI4Interconnect/_1121_ ( .A1(\AXI4Interconnect/_0743_ ), .A2(\AXI4Interconnect/_0739_ ), .A3(\AXI4Interconnect/_0744_ ), .A4(\AXI4Interconnect/_0745_ ), .ZN(\AXI4Interconnect/_0290_ ) );
INV_X1 \AXI4Interconnect/_1122_ ( .A(\AXI4Interconnect/_0141_ ), .ZN(\AXI4Interconnect/_0746_ ) );
NOR4_X1 \AXI4Interconnect/_1123_ ( .A1(\AXI4Interconnect/_0743_ ), .A2(\AXI4Interconnect/_0739_ ), .A3(\AXI4Interconnect/_0744_ ), .A4(\AXI4Interconnect/_0746_ ), .ZN(\AXI4Interconnect/_0291_ ) );
INV_X1 \AXI4Interconnect/_1124_ ( .A(\AXI4Interconnect/_0194_ ), .ZN(\AXI4Interconnect/_0747_ ) );
NOR4_X1 \AXI4Interconnect/_1125_ ( .A1(\AXI4Interconnect/_0743_ ), .A2(\AXI4Interconnect/_0739_ ), .A3(\AXI4Interconnect/_0744_ ), .A4(\AXI4Interconnect/_0747_ ), .ZN(\AXI4Interconnect/_0341_ ) );
INV_X1 \AXI4Interconnect/_1126_ ( .A(\AXI4Interconnect/_0205_ ), .ZN(\AXI4Interconnect/_0748_ ) );
NOR4_X1 \AXI4Interconnect/_1127_ ( .A1(\AXI4Interconnect/_0743_ ), .A2(\AXI4Interconnect/_0739_ ), .A3(\AXI4Interconnect/_0744_ ), .A4(\AXI4Interconnect/_0748_ ), .ZN(\AXI4Interconnect/_0352_ ) );
INV_X1 \AXI4Interconnect/_1128_ ( .A(\AXI4Interconnect/_0216_ ), .ZN(\AXI4Interconnect/_0749_ ) );
NOR4_X1 \AXI4Interconnect/_1129_ ( .A1(\AXI4Interconnect/_0743_ ), .A2(\AXI4Interconnect/_0739_ ), .A3(\AXI4Interconnect/_0744_ ), .A4(\AXI4Interconnect/_0749_ ), .ZN(\AXI4Interconnect/_0363_ ) );
INV_X1 \AXI4Interconnect/_1130_ ( .A(\AXI4Interconnect/_0219_ ), .ZN(\AXI4Interconnect/_0750_ ) );
NOR4_X1 \AXI4Interconnect/_1131_ ( .A1(\AXI4Interconnect/_0743_ ), .A2(\AXI4Interconnect/_0739_ ), .A3(\AXI4Interconnect/_0744_ ), .A4(\AXI4Interconnect/_0750_ ), .ZN(\AXI4Interconnect/_0366_ ) );
INV_X1 \AXI4Interconnect/_1132_ ( .A(\AXI4Interconnect/_0220_ ), .ZN(\AXI4Interconnect/_0751_ ) );
NOR4_X1 \AXI4Interconnect/_1133_ ( .A1(\AXI4Interconnect/_0743_ ), .A2(\AXI4Interconnect/_0739_ ), .A3(\AXI4Interconnect/_0744_ ), .A4(\AXI4Interconnect/_0751_ ), .ZN(\AXI4Interconnect/_0367_ ) );
INV_X1 \AXI4Interconnect/_1134_ ( .A(\AXI4Interconnect/_0221_ ), .ZN(\AXI4Interconnect/_0752_ ) );
NOR4_X1 \AXI4Interconnect/_1135_ ( .A1(\AXI4Interconnect/_0743_ ), .A2(\AXI4Interconnect/_0739_ ), .A3(\AXI4Interconnect/_0744_ ), .A4(\AXI4Interconnect/_0752_ ), .ZN(\AXI4Interconnect/_0368_ ) );
BUF_X4 \AXI4Interconnect/_1136_ ( .A(\AXI4Interconnect/_0712_ ), .Z(\AXI4Interconnect/_0753_ ) );
INV_X1 \AXI4Interconnect/_1137_ ( .A(\AXI4Interconnect/_0222_ ), .ZN(\AXI4Interconnect/_0754_ ) );
NOR4_X1 \AXI4Interconnect/_1138_ ( .A1(\AXI4Interconnect/_0743_ ), .A2(\AXI4Interconnect/_0753_ ), .A3(\AXI4Interconnect/_0744_ ), .A4(\AXI4Interconnect/_0754_ ), .ZN(\AXI4Interconnect/_0369_ ) );
INV_X1 \AXI4Interconnect/_1139_ ( .A(\AXI4Interconnect/_0223_ ), .ZN(\AXI4Interconnect/_0755_ ) );
NOR4_X1 \AXI4Interconnect/_1140_ ( .A1(\AXI4Interconnect/_0743_ ), .A2(\AXI4Interconnect/_0753_ ), .A3(\AXI4Interconnect/_0744_ ), .A4(\AXI4Interconnect/_0755_ ), .ZN(\AXI4Interconnect/_0370_ ) );
BUF_X4 \AXI4Interconnect/_1141_ ( .A(\AXI4Interconnect/_0742_ ), .Z(\AXI4Interconnect/_0756_ ) );
BUF_X4 \AXI4Interconnect/_1142_ ( .A(\AXI4Interconnect/_0701_ ), .Z(\AXI4Interconnect/_0757_ ) );
INV_X1 \AXI4Interconnect/_1143_ ( .A(\AXI4Interconnect/_0224_ ), .ZN(\AXI4Interconnect/_0758_ ) );
NOR4_X1 \AXI4Interconnect/_1144_ ( .A1(\AXI4Interconnect/_0756_ ), .A2(\AXI4Interconnect/_0753_ ), .A3(\AXI4Interconnect/_0757_ ), .A4(\AXI4Interconnect/_0758_ ), .ZN(\AXI4Interconnect/_0371_ ) );
INV_X1 \AXI4Interconnect/_1145_ ( .A(\AXI4Interconnect/_0225_ ), .ZN(\AXI4Interconnect/_0759_ ) );
NOR4_X1 \AXI4Interconnect/_1146_ ( .A1(\AXI4Interconnect/_0756_ ), .A2(\AXI4Interconnect/_0753_ ), .A3(\AXI4Interconnect/_0757_ ), .A4(\AXI4Interconnect/_0759_ ), .ZN(\AXI4Interconnect/_0372_ ) );
INV_X1 \AXI4Interconnect/_1147_ ( .A(\AXI4Interconnect/_0195_ ), .ZN(\AXI4Interconnect/_0760_ ) );
NOR4_X1 \AXI4Interconnect/_1148_ ( .A1(\AXI4Interconnect/_0756_ ), .A2(\AXI4Interconnect/_0753_ ), .A3(\AXI4Interconnect/_0757_ ), .A4(\AXI4Interconnect/_0760_ ), .ZN(\AXI4Interconnect/_0342_ ) );
INV_X1 \AXI4Interconnect/_1149_ ( .A(\AXI4Interconnect/_0196_ ), .ZN(\AXI4Interconnect/_0761_ ) );
NOR4_X1 \AXI4Interconnect/_1150_ ( .A1(\AXI4Interconnect/_0756_ ), .A2(\AXI4Interconnect/_0753_ ), .A3(\AXI4Interconnect/_0757_ ), .A4(\AXI4Interconnect/_0761_ ), .ZN(\AXI4Interconnect/_0343_ ) );
INV_X1 \AXI4Interconnect/_1151_ ( .A(\AXI4Interconnect/_0197_ ), .ZN(\AXI4Interconnect/_0762_ ) );
NOR4_X1 \AXI4Interconnect/_1152_ ( .A1(\AXI4Interconnect/_0756_ ), .A2(\AXI4Interconnect/_0753_ ), .A3(\AXI4Interconnect/_0757_ ), .A4(\AXI4Interconnect/_0762_ ), .ZN(\AXI4Interconnect/_0344_ ) );
INV_X1 \AXI4Interconnect/_1153_ ( .A(\AXI4Interconnect/_0198_ ), .ZN(\AXI4Interconnect/_0763_ ) );
NOR4_X1 \AXI4Interconnect/_1154_ ( .A1(\AXI4Interconnect/_0756_ ), .A2(\AXI4Interconnect/_0753_ ), .A3(\AXI4Interconnect/_0757_ ), .A4(\AXI4Interconnect/_0763_ ), .ZN(\AXI4Interconnect/_0345_ ) );
INV_X1 \AXI4Interconnect/_1155_ ( .A(\AXI4Interconnect/_0199_ ), .ZN(\AXI4Interconnect/_0764_ ) );
NOR4_X1 \AXI4Interconnect/_1156_ ( .A1(\AXI4Interconnect/_0756_ ), .A2(\AXI4Interconnect/_0753_ ), .A3(\AXI4Interconnect/_0757_ ), .A4(\AXI4Interconnect/_0764_ ), .ZN(\AXI4Interconnect/_0346_ ) );
INV_X1 \AXI4Interconnect/_1157_ ( .A(\AXI4Interconnect/_0200_ ), .ZN(\AXI4Interconnect/_0765_ ) );
NOR4_X1 \AXI4Interconnect/_1158_ ( .A1(\AXI4Interconnect/_0756_ ), .A2(\AXI4Interconnect/_0753_ ), .A3(\AXI4Interconnect/_0757_ ), .A4(\AXI4Interconnect/_0765_ ), .ZN(\AXI4Interconnect/_0347_ ) );
BUF_X4 \AXI4Interconnect/_1159_ ( .A(\AXI4Interconnect/_0712_ ), .Z(\AXI4Interconnect/_0766_ ) );
INV_X1 \AXI4Interconnect/_1160_ ( .A(\AXI4Interconnect/_0201_ ), .ZN(\AXI4Interconnect/_0767_ ) );
NOR4_X1 \AXI4Interconnect/_1161_ ( .A1(\AXI4Interconnect/_0756_ ), .A2(\AXI4Interconnect/_0766_ ), .A3(\AXI4Interconnect/_0757_ ), .A4(\AXI4Interconnect/_0767_ ), .ZN(\AXI4Interconnect/_0348_ ) );
INV_X1 \AXI4Interconnect/_1162_ ( .A(\AXI4Interconnect/_0202_ ), .ZN(\AXI4Interconnect/_0768_ ) );
NOR4_X1 \AXI4Interconnect/_1163_ ( .A1(\AXI4Interconnect/_0756_ ), .A2(\AXI4Interconnect/_0766_ ), .A3(\AXI4Interconnect/_0757_ ), .A4(\AXI4Interconnect/_0768_ ), .ZN(\AXI4Interconnect/_0349_ ) );
BUF_X4 \AXI4Interconnect/_1164_ ( .A(\AXI4Interconnect/_0742_ ), .Z(\AXI4Interconnect/_0769_ ) );
BUF_X4 \AXI4Interconnect/_1165_ ( .A(\AXI4Interconnect/_0701_ ), .Z(\AXI4Interconnect/_0770_ ) );
INV_X1 \AXI4Interconnect/_1166_ ( .A(\AXI4Interconnect/_0203_ ), .ZN(\AXI4Interconnect/_0771_ ) );
NOR4_X1 \AXI4Interconnect/_1167_ ( .A1(\AXI4Interconnect/_0769_ ), .A2(\AXI4Interconnect/_0766_ ), .A3(\AXI4Interconnect/_0770_ ), .A4(\AXI4Interconnect/_0771_ ), .ZN(\AXI4Interconnect/_0350_ ) );
INV_X1 \AXI4Interconnect/_1168_ ( .A(\AXI4Interconnect/_0204_ ), .ZN(\AXI4Interconnect/_0772_ ) );
NOR4_X1 \AXI4Interconnect/_1169_ ( .A1(\AXI4Interconnect/_0769_ ), .A2(\AXI4Interconnect/_0766_ ), .A3(\AXI4Interconnect/_0770_ ), .A4(\AXI4Interconnect/_0772_ ), .ZN(\AXI4Interconnect/_0351_ ) );
INV_X1 \AXI4Interconnect/_1170_ ( .A(\AXI4Interconnect/_0206_ ), .ZN(\AXI4Interconnect/_0773_ ) );
NOR4_X1 \AXI4Interconnect/_1171_ ( .A1(\AXI4Interconnect/_0769_ ), .A2(\AXI4Interconnect/_0766_ ), .A3(\AXI4Interconnect/_0770_ ), .A4(\AXI4Interconnect/_0773_ ), .ZN(\AXI4Interconnect/_0353_ ) );
INV_X1 \AXI4Interconnect/_1172_ ( .A(\AXI4Interconnect/_0207_ ), .ZN(\AXI4Interconnect/_0774_ ) );
NOR4_X1 \AXI4Interconnect/_1173_ ( .A1(\AXI4Interconnect/_0769_ ), .A2(\AXI4Interconnect/_0766_ ), .A3(\AXI4Interconnect/_0770_ ), .A4(\AXI4Interconnect/_0774_ ), .ZN(\AXI4Interconnect/_0354_ ) );
INV_X1 \AXI4Interconnect/_1174_ ( .A(\AXI4Interconnect/_0208_ ), .ZN(\AXI4Interconnect/_0775_ ) );
NOR4_X1 \AXI4Interconnect/_1175_ ( .A1(\AXI4Interconnect/_0769_ ), .A2(\AXI4Interconnect/_0766_ ), .A3(\AXI4Interconnect/_0770_ ), .A4(\AXI4Interconnect/_0775_ ), .ZN(\AXI4Interconnect/_0355_ ) );
INV_X1 \AXI4Interconnect/_1176_ ( .A(\AXI4Interconnect/_0209_ ), .ZN(\AXI4Interconnect/_0776_ ) );
NOR4_X1 \AXI4Interconnect/_1177_ ( .A1(\AXI4Interconnect/_0769_ ), .A2(\AXI4Interconnect/_0766_ ), .A3(\AXI4Interconnect/_0770_ ), .A4(\AXI4Interconnect/_0776_ ), .ZN(\AXI4Interconnect/_0356_ ) );
INV_X1 \AXI4Interconnect/_1178_ ( .A(\AXI4Interconnect/_0210_ ), .ZN(\AXI4Interconnect/_0777_ ) );
NOR4_X1 \AXI4Interconnect/_1179_ ( .A1(\AXI4Interconnect/_0769_ ), .A2(\AXI4Interconnect/_0766_ ), .A3(\AXI4Interconnect/_0770_ ), .A4(\AXI4Interconnect/_0777_ ), .ZN(\AXI4Interconnect/_0357_ ) );
INV_X1 \AXI4Interconnect/_1180_ ( .A(\AXI4Interconnect/_0211_ ), .ZN(\AXI4Interconnect/_0778_ ) );
NOR4_X1 \AXI4Interconnect/_1181_ ( .A1(\AXI4Interconnect/_0769_ ), .A2(\AXI4Interconnect/_0766_ ), .A3(\AXI4Interconnect/_0770_ ), .A4(\AXI4Interconnect/_0778_ ), .ZN(\AXI4Interconnect/_0358_ ) );
BUF_X4 \AXI4Interconnect/_1182_ ( .A(\AXI4Interconnect/_0712_ ), .Z(\AXI4Interconnect/_0779_ ) );
INV_X1 \AXI4Interconnect/_1183_ ( .A(\AXI4Interconnect/_0212_ ), .ZN(\AXI4Interconnect/_0780_ ) );
NOR4_X1 \AXI4Interconnect/_1184_ ( .A1(\AXI4Interconnect/_0769_ ), .A2(\AXI4Interconnect/_0779_ ), .A3(\AXI4Interconnect/_0770_ ), .A4(\AXI4Interconnect/_0780_ ), .ZN(\AXI4Interconnect/_0359_ ) );
INV_X1 \AXI4Interconnect/_1185_ ( .A(\AXI4Interconnect/_0213_ ), .ZN(\AXI4Interconnect/_0781_ ) );
NOR4_X1 \AXI4Interconnect/_1186_ ( .A1(\AXI4Interconnect/_0769_ ), .A2(\AXI4Interconnect/_0779_ ), .A3(\AXI4Interconnect/_0770_ ), .A4(\AXI4Interconnect/_0781_ ), .ZN(\AXI4Interconnect/_0360_ ) );
BUF_X4 \AXI4Interconnect/_1187_ ( .A(\AXI4Interconnect/_0742_ ), .Z(\AXI4Interconnect/_0782_ ) );
INV_X1 \AXI4Interconnect/_1188_ ( .A(\AXI4Interconnect/_0214_ ), .ZN(\AXI4Interconnect/_0783_ ) );
NOR4_X1 \AXI4Interconnect/_1189_ ( .A1(\AXI4Interconnect/_0782_ ), .A2(\AXI4Interconnect/_0779_ ), .A3(\AXI4Interconnect/_0702_ ), .A4(\AXI4Interconnect/_0783_ ), .ZN(\AXI4Interconnect/_0361_ ) );
INV_X1 \AXI4Interconnect/_1190_ ( .A(\AXI4Interconnect/_0215_ ), .ZN(\AXI4Interconnect/_0784_ ) );
NOR4_X1 \AXI4Interconnect/_1191_ ( .A1(\AXI4Interconnect/_0782_ ), .A2(\AXI4Interconnect/_0779_ ), .A3(\AXI4Interconnect/_0702_ ), .A4(\AXI4Interconnect/_0784_ ), .ZN(\AXI4Interconnect/_0362_ ) );
INV_X1 \AXI4Interconnect/_1192_ ( .A(\AXI4Interconnect/_0217_ ), .ZN(\AXI4Interconnect/_0785_ ) );
NOR4_X1 \AXI4Interconnect/_1193_ ( .A1(\AXI4Interconnect/_0782_ ), .A2(\AXI4Interconnect/_0779_ ), .A3(\AXI4Interconnect/_0702_ ), .A4(\AXI4Interconnect/_0785_ ), .ZN(\AXI4Interconnect/_0364_ ) );
INV_X1 \AXI4Interconnect/_1194_ ( .A(\AXI4Interconnect/_0218_ ), .ZN(\AXI4Interconnect/_0786_ ) );
NOR4_X1 \AXI4Interconnect/_1195_ ( .A1(\AXI4Interconnect/_0782_ ), .A2(\AXI4Interconnect/_0779_ ), .A3(\AXI4Interconnect/_0702_ ), .A4(\AXI4Interconnect/_0786_ ), .ZN(\AXI4Interconnect/_0365_ ) );
NOR2_X1 \AXI4Interconnect/_1196_ ( .A1(\AXI4Interconnect/_0611_ ), .A2(\AXI4Interconnect/_0701_ ), .ZN(\AXI4Interconnect/_0787_ ) );
INV_X1 \AXI4Interconnect/_1197_ ( .A(\AXI4Interconnect/_0787_ ), .ZN(\AXI4Interconnect/_0788_ ) );
BUF_X4 \AXI4Interconnect/_1198_ ( .A(\AXI4Interconnect/_0788_ ), .Z(\AXI4Interconnect/_0789_ ) );
OR2_X1 \AXI4Interconnect/_1199_ ( .A1(fanout_net_6 ), .A2(\AXI4Interconnect/_0010_ ), .ZN(\AXI4Interconnect/_0790_ ) );
BUF_X4 \AXI4Interconnect/_1200_ ( .A(\AXI4Interconnect/_0712_ ), .Z(\AXI4Interconnect/_0791_ ) );
OAI21_X1 \AXI4Interconnect/_1201_ ( .A(\AXI4Interconnect/_0790_ ), .B1(\AXI4Interconnect/_0791_ ), .B2(\AXI4Interconnect/_0080_ ), .ZN(\AXI4Interconnect/_0792_ ) );
NOR2_X1 \AXI4Interconnect/_1202_ ( .A1(\AXI4Interconnect/_0789_ ), .A2(\AXI4Interconnect/_0792_ ), .ZN(\AXI4Interconnect/_0233_ ) );
OR2_X1 \AXI4Interconnect/_1203_ ( .A1(fanout_net_6 ), .A2(\AXI4Interconnect/_0021_ ), .ZN(\AXI4Interconnect/_0793_ ) );
OAI21_X1 \AXI4Interconnect/_1204_ ( .A(\AXI4Interconnect/_0793_ ), .B1(\AXI4Interconnect/_0791_ ), .B2(\AXI4Interconnect/_0091_ ), .ZN(\AXI4Interconnect/_0794_ ) );
NOR2_X1 \AXI4Interconnect/_1205_ ( .A1(\AXI4Interconnect/_0789_ ), .A2(\AXI4Interconnect/_0794_ ), .ZN(\AXI4Interconnect/_0244_ ) );
AND2_X1 \AXI4Interconnect/_1206_ ( .A1(fanout_net_6 ), .A2(\AXI4Interconnect/_0102_ ), .ZN(\AXI4Interconnect/_0795_ ) );
AOI21_X1 \AXI4Interconnect/_1207_ ( .A(\AXI4Interconnect/_0795_ ), .B1(\AXI4Interconnect/_0791_ ), .B2(\AXI4Interconnect/_0032_ ), .ZN(\AXI4Interconnect/_0796_ ) );
NOR2_X1 \AXI4Interconnect/_1208_ ( .A1(\AXI4Interconnect/_0789_ ), .A2(\AXI4Interconnect/_0796_ ), .ZN(\AXI4Interconnect/_0255_ ) );
OR2_X1 \AXI4Interconnect/_1209_ ( .A1(fanout_net_6 ), .A2(\AXI4Interconnect/_0035_ ), .ZN(\AXI4Interconnect/_0797_ ) );
OAI21_X1 \AXI4Interconnect/_1210_ ( .A(\AXI4Interconnect/_0797_ ), .B1(\AXI4Interconnect/_0791_ ), .B2(\AXI4Interconnect/_0105_ ), .ZN(\AXI4Interconnect/_0798_ ) );
NOR2_X1 \AXI4Interconnect/_1211_ ( .A1(\AXI4Interconnect/_0789_ ), .A2(\AXI4Interconnect/_0798_ ), .ZN(\AXI4Interconnect/_0258_ ) );
OR2_X1 \AXI4Interconnect/_1212_ ( .A1(fanout_net_6 ), .A2(\AXI4Interconnect/_0036_ ), .ZN(\AXI4Interconnect/_0799_ ) );
OAI21_X1 \AXI4Interconnect/_1213_ ( .A(\AXI4Interconnect/_0799_ ), .B1(\AXI4Interconnect/_0791_ ), .B2(\AXI4Interconnect/_0106_ ), .ZN(\AXI4Interconnect/_0800_ ) );
NOR2_X1 \AXI4Interconnect/_1214_ ( .A1(\AXI4Interconnect/_0789_ ), .A2(\AXI4Interconnect/_0800_ ), .ZN(\AXI4Interconnect/_0259_ ) );
AND2_X1 \AXI4Interconnect/_1215_ ( .A1(fanout_net_6 ), .A2(\AXI4Interconnect/_0107_ ), .ZN(\AXI4Interconnect/_0801_ ) );
AOI21_X1 \AXI4Interconnect/_1216_ ( .A(\AXI4Interconnect/_0801_ ), .B1(\AXI4Interconnect/_0791_ ), .B2(\AXI4Interconnect/_0037_ ), .ZN(\AXI4Interconnect/_0802_ ) );
NOR2_X1 \AXI4Interconnect/_1217_ ( .A1(\AXI4Interconnect/_0789_ ), .A2(\AXI4Interconnect/_0802_ ), .ZN(\AXI4Interconnect/_0260_ ) );
AND2_X1 \AXI4Interconnect/_1218_ ( .A1(fanout_net_6 ), .A2(\AXI4Interconnect/_0108_ ), .ZN(\AXI4Interconnect/_0803_ ) );
AOI21_X1 \AXI4Interconnect/_1219_ ( .A(\AXI4Interconnect/_0803_ ), .B1(\AXI4Interconnect/_0791_ ), .B2(\AXI4Interconnect/_0038_ ), .ZN(\AXI4Interconnect/_0804_ ) );
NOR2_X1 \AXI4Interconnect/_1220_ ( .A1(\AXI4Interconnect/_0789_ ), .A2(\AXI4Interconnect/_0804_ ), .ZN(\AXI4Interconnect/_0261_ ) );
AND2_X1 \AXI4Interconnect/_1221_ ( .A1(\AXI4Interconnect/_0712_ ), .A2(\AXI4Interconnect/_0039_ ), .ZN(\AXI4Interconnect/_0805_ ) );
AOI21_X1 \AXI4Interconnect/_1222_ ( .A(\AXI4Interconnect/_0805_ ), .B1(fanout_net_6 ), .B2(\AXI4Interconnect/_0109_ ), .ZN(\AXI4Interconnect/_0806_ ) );
BUF_X4 \AXI4Interconnect/_1223_ ( .A(\AXI4Interconnect/_0788_ ), .Z(\AXI4Interconnect/_0807_ ) );
NOR2_X1 \AXI4Interconnect/_1224_ ( .A1(\AXI4Interconnect/_0806_ ), .A2(\AXI4Interconnect/_0807_ ), .ZN(\AXI4Interconnect/_0262_ ) );
OR2_X1 \AXI4Interconnect/_1225_ ( .A1(\AXI4Interconnect/_0712_ ), .A2(\AXI4Interconnect/_0110_ ), .ZN(\AXI4Interconnect/_0808_ ) );
OAI21_X1 \AXI4Interconnect/_1226_ ( .A(\AXI4Interconnect/_0808_ ), .B1(fanout_net_6 ), .B2(\AXI4Interconnect/_0040_ ), .ZN(\AXI4Interconnect/_0809_ ) );
NOR2_X1 \AXI4Interconnect/_1227_ ( .A1(\AXI4Interconnect/_0809_ ), .A2(\AXI4Interconnect/_0807_ ), .ZN(\AXI4Interconnect/_0263_ ) );
AND2_X1 \AXI4Interconnect/_1228_ ( .A1(\AXI4Interconnect/_0698_ ), .A2(\AXI4Interconnect/_0041_ ), .ZN(\AXI4Interconnect/_0810_ ) );
AOI21_X1 \AXI4Interconnect/_1229_ ( .A(\AXI4Interconnect/_0810_ ), .B1(fanout_net_6 ), .B2(\AXI4Interconnect/_0111_ ), .ZN(\AXI4Interconnect/_0811_ ) );
NOR2_X1 \AXI4Interconnect/_1230_ ( .A1(\AXI4Interconnect/_0811_ ), .A2(\AXI4Interconnect/_0807_ ), .ZN(\AXI4Interconnect/_0264_ ) );
AND2_X1 \AXI4Interconnect/_1231_ ( .A1(fanout_net_6 ), .A2(\AXI4Interconnect/_0081_ ), .ZN(\AXI4Interconnect/_0812_ ) );
AOI21_X1 \AXI4Interconnect/_1232_ ( .A(\AXI4Interconnect/_0812_ ), .B1(\AXI4Interconnect/_0791_ ), .B2(\AXI4Interconnect/_0011_ ), .ZN(\AXI4Interconnect/_0813_ ) );
NOR2_X1 \AXI4Interconnect/_1233_ ( .A1(\AXI4Interconnect/_0789_ ), .A2(\AXI4Interconnect/_0813_ ), .ZN(\AXI4Interconnect/_0234_ ) );
AND2_X1 \AXI4Interconnect/_1234_ ( .A1(fanout_net_6 ), .A2(\AXI4Interconnect/_0082_ ), .ZN(\AXI4Interconnect/_0814_ ) );
AOI21_X1 \AXI4Interconnect/_1235_ ( .A(\AXI4Interconnect/_0814_ ), .B1(\AXI4Interconnect/_0791_ ), .B2(\AXI4Interconnect/_0012_ ), .ZN(\AXI4Interconnect/_0815_ ) );
NOR2_X1 \AXI4Interconnect/_1236_ ( .A1(\AXI4Interconnect/_0789_ ), .A2(\AXI4Interconnect/_0815_ ), .ZN(\AXI4Interconnect/_0235_ ) );
AND2_X1 \AXI4Interconnect/_1237_ ( .A1(\AXI4Interconnect/_0698_ ), .A2(\AXI4Interconnect/_0013_ ), .ZN(\AXI4Interconnect/_0816_ ) );
AOI21_X1 \AXI4Interconnect/_1238_ ( .A(\AXI4Interconnect/_0816_ ), .B1(fanout_net_6 ), .B2(\AXI4Interconnect/_0083_ ), .ZN(\AXI4Interconnect/_0817_ ) );
NOR2_X1 \AXI4Interconnect/_1239_ ( .A1(\AXI4Interconnect/_0817_ ), .A2(\AXI4Interconnect/_0807_ ), .ZN(\AXI4Interconnect/_0236_ ) );
AND2_X1 \AXI4Interconnect/_1240_ ( .A1(\AXI4Interconnect/_0698_ ), .A2(\AXI4Interconnect/_0014_ ), .ZN(\AXI4Interconnect/_0818_ ) );
AOI21_X1 \AXI4Interconnect/_1241_ ( .A(\AXI4Interconnect/_0818_ ), .B1(fanout_net_6 ), .B2(\AXI4Interconnect/_0084_ ), .ZN(\AXI4Interconnect/_0819_ ) );
NOR2_X1 \AXI4Interconnect/_1242_ ( .A1(\AXI4Interconnect/_0819_ ), .A2(\AXI4Interconnect/_0807_ ), .ZN(\AXI4Interconnect/_0237_ ) );
OR2_X1 \AXI4Interconnect/_1243_ ( .A1(fanout_net_6 ), .A2(\AXI4Interconnect/_0015_ ), .ZN(\AXI4Interconnect/_0820_ ) );
OAI21_X1 \AXI4Interconnect/_1244_ ( .A(\AXI4Interconnect/_0820_ ), .B1(\AXI4Interconnect/_0699_ ), .B2(\AXI4Interconnect/_0085_ ), .ZN(\AXI4Interconnect/_0821_ ) );
NOR2_X1 \AXI4Interconnect/_1245_ ( .A1(\AXI4Interconnect/_0789_ ), .A2(\AXI4Interconnect/_0821_ ), .ZN(\AXI4Interconnect/_0238_ ) );
BUF_X4 \AXI4Interconnect/_1246_ ( .A(\AXI4Interconnect/_0788_ ), .Z(\AXI4Interconnect/_0822_ ) );
OR2_X1 \AXI4Interconnect/_1247_ ( .A1(fanout_net_6 ), .A2(\AXI4Interconnect/_0016_ ), .ZN(\AXI4Interconnect/_0823_ ) );
OAI21_X1 \AXI4Interconnect/_1248_ ( .A(\AXI4Interconnect/_0823_ ), .B1(\AXI4Interconnect/_0699_ ), .B2(\AXI4Interconnect/_0086_ ), .ZN(\AXI4Interconnect/_0824_ ) );
NOR2_X1 \AXI4Interconnect/_1249_ ( .A1(\AXI4Interconnect/_0822_ ), .A2(\AXI4Interconnect/_0824_ ), .ZN(\AXI4Interconnect/_0239_ ) );
OR2_X1 \AXI4Interconnect/_1250_ ( .A1(fanout_net_6 ), .A2(\AXI4Interconnect/_0017_ ), .ZN(\AXI4Interconnect/_0825_ ) );
OAI21_X1 \AXI4Interconnect/_1251_ ( .A(\AXI4Interconnect/_0825_ ), .B1(\AXI4Interconnect/_0699_ ), .B2(\AXI4Interconnect/_0087_ ), .ZN(\AXI4Interconnect/_0826_ ) );
NOR2_X1 \AXI4Interconnect/_1252_ ( .A1(\AXI4Interconnect/_0822_ ), .A2(\AXI4Interconnect/_0826_ ), .ZN(\AXI4Interconnect/_0240_ ) );
OR2_X1 \AXI4Interconnect/_1253_ ( .A1(fanout_net_6 ), .A2(\AXI4Interconnect/_0018_ ), .ZN(\AXI4Interconnect/_0827_ ) );
OAI21_X1 \AXI4Interconnect/_1254_ ( .A(\AXI4Interconnect/_0827_ ), .B1(\AXI4Interconnect/_0699_ ), .B2(\AXI4Interconnect/_0088_ ), .ZN(\AXI4Interconnect/_0828_ ) );
NOR2_X1 \AXI4Interconnect/_1255_ ( .A1(\AXI4Interconnect/_0822_ ), .A2(\AXI4Interconnect/_0828_ ), .ZN(\AXI4Interconnect/_0241_ ) );
OR2_X1 \AXI4Interconnect/_1256_ ( .A1(fanout_net_6 ), .A2(\AXI4Interconnect/_0019_ ), .ZN(\AXI4Interconnect/_0829_ ) );
OAI21_X1 \AXI4Interconnect/_1257_ ( .A(\AXI4Interconnect/_0829_ ), .B1(\AXI4Interconnect/_0699_ ), .B2(\AXI4Interconnect/_0089_ ), .ZN(\AXI4Interconnect/_0830_ ) );
NOR2_X1 \AXI4Interconnect/_1258_ ( .A1(\AXI4Interconnect/_0822_ ), .A2(\AXI4Interconnect/_0830_ ), .ZN(\AXI4Interconnect/_0242_ ) );
AND2_X1 \AXI4Interconnect/_1259_ ( .A1(\AXI4Interconnect/_0698_ ), .A2(\AXI4Interconnect/_0020_ ), .ZN(\AXI4Interconnect/_0831_ ) );
AOI21_X1 \AXI4Interconnect/_1260_ ( .A(\AXI4Interconnect/_0831_ ), .B1(fanout_net_6 ), .B2(\AXI4Interconnect/_0090_ ), .ZN(\AXI4Interconnect/_0832_ ) );
NOR2_X1 \AXI4Interconnect/_1261_ ( .A1(\AXI4Interconnect/_0832_ ), .A2(\AXI4Interconnect/_0807_ ), .ZN(\AXI4Interconnect/_0243_ ) );
OR2_X1 \AXI4Interconnect/_1262_ ( .A1(fanout_net_6 ), .A2(\AXI4Interconnect/_0022_ ), .ZN(\AXI4Interconnect/_0833_ ) );
OAI21_X1 \AXI4Interconnect/_1263_ ( .A(\AXI4Interconnect/_0833_ ), .B1(\AXI4Interconnect/_0699_ ), .B2(\AXI4Interconnect/_0092_ ), .ZN(\AXI4Interconnect/_0834_ ) );
NOR2_X1 \AXI4Interconnect/_1264_ ( .A1(\AXI4Interconnect/_0822_ ), .A2(\AXI4Interconnect/_0834_ ), .ZN(\AXI4Interconnect/_0245_ ) );
AND2_X1 \AXI4Interconnect/_1265_ ( .A1(\AXI4Interconnect/_0698_ ), .A2(\AXI4Interconnect/_0023_ ), .ZN(\AXI4Interconnect/_0835_ ) );
AOI21_X1 \AXI4Interconnect/_1266_ ( .A(\AXI4Interconnect/_0835_ ), .B1(fanout_net_6 ), .B2(\AXI4Interconnect/_0093_ ), .ZN(\AXI4Interconnect/_0836_ ) );
NOR2_X1 \AXI4Interconnect/_1267_ ( .A1(\AXI4Interconnect/_0836_ ), .A2(\AXI4Interconnect/_0807_ ), .ZN(\AXI4Interconnect/_0246_ ) );
AND2_X1 \AXI4Interconnect/_1268_ ( .A1(\AXI4Interconnect/_0698_ ), .A2(\AXI4Interconnect/_0024_ ), .ZN(\AXI4Interconnect/_0837_ ) );
AOI21_X1 \AXI4Interconnect/_1269_ ( .A(\AXI4Interconnect/_0837_ ), .B1(fanout_net_6 ), .B2(\AXI4Interconnect/_0094_ ), .ZN(\AXI4Interconnect/_0838_ ) );
NOR2_X1 \AXI4Interconnect/_1270_ ( .A1(\AXI4Interconnect/_0838_ ), .A2(\AXI4Interconnect/_0788_ ), .ZN(\AXI4Interconnect/_0247_ ) );
OR2_X1 \AXI4Interconnect/_1271_ ( .A1(\AXI4Interconnect/_0712_ ), .A2(\AXI4Interconnect/_0095_ ), .ZN(\AXI4Interconnect/_0839_ ) );
OAI21_X1 \AXI4Interconnect/_1272_ ( .A(\AXI4Interconnect/_0839_ ), .B1(fanout_net_6 ), .B2(\AXI4Interconnect/_0025_ ), .ZN(\AXI4Interconnect/_0840_ ) );
NOR2_X1 \AXI4Interconnect/_1273_ ( .A1(\AXI4Interconnect/_0840_ ), .A2(\AXI4Interconnect/_0788_ ), .ZN(\AXI4Interconnect/_0248_ ) );
AND2_X1 \AXI4Interconnect/_1274_ ( .A1(\AXI4Interconnect/_0698_ ), .A2(\AXI4Interconnect/_0026_ ), .ZN(\AXI4Interconnect/_0841_ ) );
AOI21_X1 \AXI4Interconnect/_1275_ ( .A(\AXI4Interconnect/_0841_ ), .B1(fanout_net_6 ), .B2(\AXI4Interconnect/_0096_ ), .ZN(\AXI4Interconnect/_0842_ ) );
NOR2_X1 \AXI4Interconnect/_1276_ ( .A1(\AXI4Interconnect/_0842_ ), .A2(\AXI4Interconnect/_0788_ ), .ZN(\AXI4Interconnect/_0249_ ) );
INV_X1 \AXI4Interconnect/_1277_ ( .A(\AXI4Interconnect/_0027_ ), .ZN(\AXI4Interconnect/_0843_ ) );
INV_X1 \AXI4Interconnect/_1278_ ( .A(\AXI4Interconnect/_0097_ ), .ZN(\AXI4Interconnect/_0844_ ) );
MUX2_X1 \AXI4Interconnect/_1279_ ( .A(\AXI4Interconnect/_0843_ ), .B(\AXI4Interconnect/_0844_ ), .S(fanout_net_6 ), .Z(\AXI4Interconnect/_0845_ ) );
NOR2_X1 \AXI4Interconnect/_1280_ ( .A1(\AXI4Interconnect/_0822_ ), .A2(\AXI4Interconnect/_0845_ ), .ZN(\AXI4Interconnect/_0250_ ) );
INV_X1 \AXI4Interconnect/_1281_ ( .A(\AXI4Interconnect/_0028_ ), .ZN(\AXI4Interconnect/_0846_ ) );
INV_X1 \AXI4Interconnect/_1282_ ( .A(\AXI4Interconnect/_0098_ ), .ZN(\AXI4Interconnect/_0847_ ) );
MUX2_X1 \AXI4Interconnect/_1283_ ( .A(\AXI4Interconnect/_0846_ ), .B(\AXI4Interconnect/_0847_ ), .S(fanout_net_6 ), .Z(\AXI4Interconnect/_0848_ ) );
NOR2_X1 \AXI4Interconnect/_1284_ ( .A1(\AXI4Interconnect/_0822_ ), .A2(\AXI4Interconnect/_0848_ ), .ZN(\AXI4Interconnect/_0251_ ) );
INV_X1 \AXI4Interconnect/_1285_ ( .A(\AXI4Interconnect/_0029_ ), .ZN(\AXI4Interconnect/_0849_ ) );
INV_X1 \AXI4Interconnect/_1286_ ( .A(\AXI4Interconnect/_0099_ ), .ZN(\AXI4Interconnect/_0850_ ) );
MUX2_X1 \AXI4Interconnect/_1287_ ( .A(\AXI4Interconnect/_0849_ ), .B(\AXI4Interconnect/_0850_ ), .S(fanout_net_6 ), .Z(\AXI4Interconnect/_0851_ ) );
NOR2_X1 \AXI4Interconnect/_1288_ ( .A1(\AXI4Interconnect/_0822_ ), .A2(\AXI4Interconnect/_0851_ ), .ZN(\AXI4Interconnect/_0252_ ) );
OR2_X1 \AXI4Interconnect/_1289_ ( .A1(fanout_net_6 ), .A2(\AXI4Interconnect/_0030_ ), .ZN(\AXI4Interconnect/_0852_ ) );
OAI21_X1 \AXI4Interconnect/_1290_ ( .A(\AXI4Interconnect/_0852_ ), .B1(\AXI4Interconnect/_0699_ ), .B2(\AXI4Interconnect/_0100_ ), .ZN(\AXI4Interconnect/_0853_ ) );
NOR2_X1 \AXI4Interconnect/_1291_ ( .A1(\AXI4Interconnect/_0822_ ), .A2(\AXI4Interconnect/_0853_ ), .ZN(\AXI4Interconnect/_0253_ ) );
OR2_X1 \AXI4Interconnect/_1292_ ( .A1(\AXI4Interconnect/_0871_ ), .A2(\AXI4Interconnect/_0031_ ), .ZN(\AXI4Interconnect/_0854_ ) );
OAI21_X1 \AXI4Interconnect/_1293_ ( .A(\AXI4Interconnect/_0854_ ), .B1(\AXI4Interconnect/_0699_ ), .B2(\AXI4Interconnect/_0101_ ), .ZN(\AXI4Interconnect/_0855_ ) );
NOR2_X1 \AXI4Interconnect/_1294_ ( .A1(\AXI4Interconnect/_0822_ ), .A2(\AXI4Interconnect/_0855_ ), .ZN(\AXI4Interconnect/_0254_ ) );
OR2_X1 \AXI4Interconnect/_1295_ ( .A1(\AXI4Interconnect/_0871_ ), .A2(\AXI4Interconnect/_0033_ ), .ZN(\AXI4Interconnect/_0856_ ) );
OAI21_X1 \AXI4Interconnect/_1296_ ( .A(\AXI4Interconnect/_0856_ ), .B1(\AXI4Interconnect/_0699_ ), .B2(\AXI4Interconnect/_0103_ ), .ZN(\AXI4Interconnect/_0857_ ) );
NOR2_X1 \AXI4Interconnect/_1297_ ( .A1(\AXI4Interconnect/_0807_ ), .A2(\AXI4Interconnect/_0857_ ), .ZN(\AXI4Interconnect/_0256_ ) );
AND2_X1 \AXI4Interconnect/_1298_ ( .A1(\AXI4Interconnect/_0871_ ), .A2(\AXI4Interconnect/_0104_ ), .ZN(\AXI4Interconnect/_0858_ ) );
AOI21_X1 \AXI4Interconnect/_1299_ ( .A(\AXI4Interconnect/_0858_ ), .B1(\AXI4Interconnect/_0791_ ), .B2(\AXI4Interconnect/_0034_ ), .ZN(\AXI4Interconnect/_0859_ ) );
NOR2_X1 \AXI4Interconnect/_1300_ ( .A1(\AXI4Interconnect/_0807_ ), .A2(\AXI4Interconnect/_0859_ ), .ZN(\AXI4Interconnect/_0257_ ) );
NOR2_X1 \AXI4Interconnect/_1301_ ( .A1(\AXI4Interconnect/_0611_ ), .A2(\AXI4Interconnect/_0607_ ), .ZN(\AXI4Interconnect/_0002_ ) );
CLKBUF_X2 \AXI4Interconnect/_1302_ ( .A(\AXI4Interconnect/_0612_ ), .Z(\AXI4Interconnect/_0860_ ) );
AND2_X1 \AXI4Interconnect/_1303_ ( .A1(\AXI4Interconnect/_0002_ ), .A2(\AXI4Interconnect/_0860_ ), .ZN(\AXI4Interconnect/_0003_ ) );
BUF_X4 \AXI4Interconnect/_1304_ ( .A(\AXI4Interconnect/_0622_ ), .Z(\AXI4Interconnect/_0861_ ) );
NOR4_X1 \AXI4Interconnect/_1305_ ( .A1(\AXI4Interconnect/_0782_ ), .A2(\AXI4Interconnect/_0861_ ), .A3(\AXI4Interconnect/_0704_ ), .A4(fanout_net_3 ), .ZN(\AXI4Interconnect/_0412_ ) );
NOR4_X1 \AXI4Interconnect/_1306_ ( .A1(\AXI4Interconnect/_0782_ ), .A2(\AXI4Interconnect/_0861_ ), .A3(\AXI4Interconnect/_0705_ ), .A4(fanout_net_3 ), .ZN(\AXI4Interconnect/_0423_ ) );
NOR4_X1 \AXI4Interconnect/_1307_ ( .A1(\AXI4Interconnect/_0782_ ), .A2(\AXI4Interconnect/_0861_ ), .A3(\AXI4Interconnect/_0706_ ), .A4(fanout_net_3 ), .ZN(\AXI4Interconnect/_0434_ ) );
NOR4_X1 \AXI4Interconnect/_1308_ ( .A1(\AXI4Interconnect/_0782_ ), .A2(\AXI4Interconnect/_0861_ ), .A3(\AXI4Interconnect/_0707_ ), .A4(fanout_net_3 ), .ZN(\AXI4Interconnect/_0437_ ) );
NOR4_X1 \AXI4Interconnect/_1309_ ( .A1(\AXI4Interconnect/_0782_ ), .A2(\AXI4Interconnect/_0861_ ), .A3(\AXI4Interconnect/_0708_ ), .A4(fanout_net_3 ), .ZN(\AXI4Interconnect/_0438_ ) );
NOR4_X1 \AXI4Interconnect/_1310_ ( .A1(\AXI4Interconnect/_0782_ ), .A2(\AXI4Interconnect/_0861_ ), .A3(\AXI4Interconnect/_0709_ ), .A4(fanout_net_3 ), .ZN(\AXI4Interconnect/_0439_ ) );
BUF_X4 \AXI4Interconnect/_1311_ ( .A(\AXI4Interconnect/_0742_ ), .Z(\AXI4Interconnect/_0862_ ) );
NOR4_X1 \AXI4Interconnect/_1312_ ( .A1(\AXI4Interconnect/_0862_ ), .A2(\AXI4Interconnect/_0861_ ), .A3(\AXI4Interconnect/_0710_ ), .A4(fanout_net_3 ), .ZN(\AXI4Interconnect/_0440_ ) );
NOR4_X1 \AXI4Interconnect/_1313_ ( .A1(\AXI4Interconnect/_0862_ ), .A2(\AXI4Interconnect/_0861_ ), .A3(\AXI4Interconnect/_0711_ ), .A4(fanout_net_3 ), .ZN(\AXI4Interconnect/_0441_ ) );
NOR4_X1 \AXI4Interconnect/_1314_ ( .A1(\AXI4Interconnect/_0862_ ), .A2(\AXI4Interconnect/_0861_ ), .A3(\AXI4Interconnect/_0714_ ), .A4(fanout_net_3 ), .ZN(\AXI4Interconnect/_0442_ ) );
BUF_X4 \AXI4Interconnect/_1315_ ( .A(\AXI4Interconnect/_0608_ ), .Z(\AXI4Interconnect/_0863_ ) );
NOR4_X1 \AXI4Interconnect/_1316_ ( .A1(\AXI4Interconnect/_0862_ ), .A2(\AXI4Interconnect/_0863_ ), .A3(\AXI4Interconnect/_0715_ ), .A4(fanout_net_3 ), .ZN(\AXI4Interconnect/_0443_ ) );
NOR4_X1 \AXI4Interconnect/_1317_ ( .A1(\AXI4Interconnect/_0862_ ), .A2(\AXI4Interconnect/_0863_ ), .A3(\AXI4Interconnect/_0718_ ), .A4(fanout_net_3 ), .ZN(\AXI4Interconnect/_0413_ ) );
NOR4_X1 \AXI4Interconnect/_1318_ ( .A1(\AXI4Interconnect/_0862_ ), .A2(\AXI4Interconnect/_0863_ ), .A3(\AXI4Interconnect/_0719_ ), .A4(fanout_net_3 ), .ZN(\AXI4Interconnect/_0414_ ) );
NOR4_X1 \AXI4Interconnect/_1319_ ( .A1(\AXI4Interconnect/_0862_ ), .A2(\AXI4Interconnect/_0863_ ), .A3(\AXI4Interconnect/_0720_ ), .A4(fanout_net_3 ), .ZN(\AXI4Interconnect/_0415_ ) );
NOR4_X1 \AXI4Interconnect/_1320_ ( .A1(\AXI4Interconnect/_0862_ ), .A2(\AXI4Interconnect/_0863_ ), .A3(\AXI4Interconnect/_0721_ ), .A4(fanout_net_3 ), .ZN(\AXI4Interconnect/_0416_ ) );
NOR4_X1 \AXI4Interconnect/_1321_ ( .A1(\AXI4Interconnect/_0862_ ), .A2(\AXI4Interconnect/_0863_ ), .A3(\AXI4Interconnect/_0722_ ), .A4(fanout_net_3 ), .ZN(\AXI4Interconnect/_0417_ ) );
NOR4_X1 \AXI4Interconnect/_1322_ ( .A1(\AXI4Interconnect/_0862_ ), .A2(\AXI4Interconnect/_0863_ ), .A3(\AXI4Interconnect/_0723_ ), .A4(fanout_net_3 ), .ZN(\AXI4Interconnect/_0418_ ) );
BUF_X4 \AXI4Interconnect/_1323_ ( .A(\AXI4Interconnect/_0742_ ), .Z(\AXI4Interconnect/_0864_ ) );
NOR4_X1 \AXI4Interconnect/_1324_ ( .A1(\AXI4Interconnect/_0864_ ), .A2(\AXI4Interconnect/_0863_ ), .A3(\AXI4Interconnect/_0724_ ), .A4(fanout_net_3 ), .ZN(\AXI4Interconnect/_0419_ ) );
NOR4_X1 \AXI4Interconnect/_1325_ ( .A1(\AXI4Interconnect/_0864_ ), .A2(\AXI4Interconnect/_0863_ ), .A3(\AXI4Interconnect/_0725_ ), .A4(fanout_net_3 ), .ZN(\AXI4Interconnect/_0420_ ) );
NOR4_X1 \AXI4Interconnect/_1326_ ( .A1(\AXI4Interconnect/_0864_ ), .A2(\AXI4Interconnect/_0863_ ), .A3(\AXI4Interconnect/_0727_ ), .A4(fanout_net_3 ), .ZN(\AXI4Interconnect/_0421_ ) );
BUF_X4 \AXI4Interconnect/_1327_ ( .A(\AXI4Interconnect/_0608_ ), .Z(\AXI4Interconnect/_0865_ ) );
NOR4_X1 \AXI4Interconnect/_1328_ ( .A1(\AXI4Interconnect/_0864_ ), .A2(\AXI4Interconnect/_0865_ ), .A3(\AXI4Interconnect/_0728_ ), .A4(fanout_net_3 ), .ZN(\AXI4Interconnect/_0422_ ) );
NOR4_X1 \AXI4Interconnect/_1329_ ( .A1(\AXI4Interconnect/_0864_ ), .A2(\AXI4Interconnect/_0865_ ), .A3(\AXI4Interconnect/_0731_ ), .A4(fanout_net_3 ), .ZN(\AXI4Interconnect/_0424_ ) );
NOR4_X1 \AXI4Interconnect/_1330_ ( .A1(\AXI4Interconnect/_0864_ ), .A2(\AXI4Interconnect/_0865_ ), .A3(\AXI4Interconnect/_0732_ ), .A4(fanout_net_3 ), .ZN(\AXI4Interconnect/_0425_ ) );
NOR4_X1 \AXI4Interconnect/_1331_ ( .A1(\AXI4Interconnect/_0864_ ), .A2(\AXI4Interconnect/_0865_ ), .A3(\AXI4Interconnect/_0733_ ), .A4(fanout_net_3 ), .ZN(\AXI4Interconnect/_0426_ ) );
NOR4_X1 \AXI4Interconnect/_1332_ ( .A1(\AXI4Interconnect/_0864_ ), .A2(\AXI4Interconnect/_0865_ ), .A3(\AXI4Interconnect/_0734_ ), .A4(fanout_net_3 ), .ZN(\AXI4Interconnect/_0427_ ) );
NOR4_X1 \AXI4Interconnect/_1333_ ( .A1(\AXI4Interconnect/_0864_ ), .A2(\AXI4Interconnect/_0865_ ), .A3(\AXI4Interconnect/_0735_ ), .A4(fanout_net_3 ), .ZN(\AXI4Interconnect/_0428_ ) );
NOR4_X1 \AXI4Interconnect/_1334_ ( .A1(\AXI4Interconnect/_0864_ ), .A2(\AXI4Interconnect/_0865_ ), .A3(\AXI4Interconnect/_0736_ ), .A4(fanout_net_3 ), .ZN(\AXI4Interconnect/_0429_ ) );
BUF_X4 \AXI4Interconnect/_1335_ ( .A(\AXI4Interconnect/_0742_ ), .Z(\AXI4Interconnect/_0866_ ) );
NOR4_X1 \AXI4Interconnect/_1336_ ( .A1(\AXI4Interconnect/_0866_ ), .A2(\AXI4Interconnect/_0865_ ), .A3(\AXI4Interconnect/_0737_ ), .A4(fanout_net_3 ), .ZN(\AXI4Interconnect/_0430_ ) );
NOR4_X1 \AXI4Interconnect/_1337_ ( .A1(\AXI4Interconnect/_0866_ ), .A2(\AXI4Interconnect/_0865_ ), .A3(\AXI4Interconnect/_0738_ ), .A4(fanout_net_3 ), .ZN(\AXI4Interconnect/_0431_ ) );
NOR4_X1 \AXI4Interconnect/_1338_ ( .A1(\AXI4Interconnect/_0866_ ), .A2(\AXI4Interconnect/_0865_ ), .A3(\AXI4Interconnect/_0740_ ), .A4(fanout_net_3 ), .ZN(\AXI4Interconnect/_0432_ ) );
BUF_X4 \AXI4Interconnect/_1339_ ( .A(\AXI4Interconnect/_0622_ ), .Z(\AXI4Interconnect/_0867_ ) );
NOR4_X1 \AXI4Interconnect/_1340_ ( .A1(\AXI4Interconnect/_0866_ ), .A2(\AXI4Interconnect/_0867_ ), .A3(\AXI4Interconnect/_0741_ ), .A4(fanout_net_4 ), .ZN(\AXI4Interconnect/_0433_ ) );
NOR4_X1 \AXI4Interconnect/_1341_ ( .A1(\AXI4Interconnect/_0866_ ), .A2(\AXI4Interconnect/_0867_ ), .A3(\AXI4Interconnect/_0745_ ), .A4(fanout_net_4 ), .ZN(\AXI4Interconnect/_0435_ ) );
NOR4_X1 \AXI4Interconnect/_1342_ ( .A1(\AXI4Interconnect/_0866_ ), .A2(\AXI4Interconnect/_0867_ ), .A3(\AXI4Interconnect/_0746_ ), .A4(fanout_net_4 ), .ZN(\AXI4Interconnect/_0436_ ) );
NOR4_X1 \AXI4Interconnect/_1343_ ( .A1(\AXI4Interconnect/_0866_ ), .A2(\AXI4Interconnect/_0867_ ), .A3(\AXI4Interconnect/_0747_ ), .A4(fanout_net_4 ), .ZN(\AXI4Interconnect/_0489_ ) );
NOR4_X1 \AXI4Interconnect/_1344_ ( .A1(\AXI4Interconnect/_0866_ ), .A2(\AXI4Interconnect/_0867_ ), .A3(\AXI4Interconnect/_0748_ ), .A4(fanout_net_4 ), .ZN(\AXI4Interconnect/_0500_ ) );
NOR4_X1 \AXI4Interconnect/_1345_ ( .A1(\AXI4Interconnect/_0866_ ), .A2(\AXI4Interconnect/_0867_ ), .A3(\AXI4Interconnect/_0749_ ), .A4(fanout_net_4 ), .ZN(\AXI4Interconnect/_0511_ ) );
NOR4_X1 \AXI4Interconnect/_1346_ ( .A1(\AXI4Interconnect/_0866_ ), .A2(\AXI4Interconnect/_0867_ ), .A3(\AXI4Interconnect/_0750_ ), .A4(fanout_net_4 ), .ZN(\AXI4Interconnect/_0514_ ) );
BUF_X4 \AXI4Interconnect/_1347_ ( .A(\AXI4Interconnect/_0742_ ), .Z(\AXI4Interconnect/_0868_ ) );
NOR4_X1 \AXI4Interconnect/_1348_ ( .A1(\AXI4Interconnect/_0868_ ), .A2(\AXI4Interconnect/_0867_ ), .A3(\AXI4Interconnect/_0751_ ), .A4(fanout_net_4 ), .ZN(\AXI4Interconnect/_0515_ ) );
NOR4_X1 \AXI4Interconnect/_1349_ ( .A1(\AXI4Interconnect/_0868_ ), .A2(\AXI4Interconnect/_0867_ ), .A3(\AXI4Interconnect/_0752_ ), .A4(fanout_net_4 ), .ZN(\AXI4Interconnect/_0516_ ) );
NOR4_X1 \AXI4Interconnect/_1350_ ( .A1(\AXI4Interconnect/_0868_ ), .A2(\AXI4Interconnect/_0867_ ), .A3(\AXI4Interconnect/_0754_ ), .A4(fanout_net_4 ), .ZN(\AXI4Interconnect/_0517_ ) );
BUF_X4 \AXI4Interconnect/_1351_ ( .A(\AXI4Interconnect/_0622_ ), .Z(\AXI4Interconnect/_0528_ ) );
NOR4_X1 \AXI4Interconnect/_1352_ ( .A1(\AXI4Interconnect/_0868_ ), .A2(\AXI4Interconnect/_0528_ ), .A3(\AXI4Interconnect/_0755_ ), .A4(fanout_net_4 ), .ZN(\AXI4Interconnect/_0518_ ) );
NOR4_X1 \AXI4Interconnect/_1353_ ( .A1(\AXI4Interconnect/_0868_ ), .A2(\AXI4Interconnect/_0528_ ), .A3(\AXI4Interconnect/_0758_ ), .A4(fanout_net_4 ), .ZN(\AXI4Interconnect/_0519_ ) );
NOR4_X1 \AXI4Interconnect/_1354_ ( .A1(\AXI4Interconnect/_0868_ ), .A2(\AXI4Interconnect/_0528_ ), .A3(\AXI4Interconnect/_0759_ ), .A4(fanout_net_4 ), .ZN(\AXI4Interconnect/_0520_ ) );
NOR4_X1 \AXI4Interconnect/_1355_ ( .A1(\AXI4Interconnect/_0868_ ), .A2(\AXI4Interconnect/_0528_ ), .A3(\AXI4Interconnect/_0760_ ), .A4(fanout_net_4 ), .ZN(\AXI4Interconnect/_0490_ ) );
NOR4_X1 \AXI4Interconnect/_1356_ ( .A1(\AXI4Interconnect/_0868_ ), .A2(\AXI4Interconnect/_0528_ ), .A3(\AXI4Interconnect/_0761_ ), .A4(fanout_net_4 ), .ZN(\AXI4Interconnect/_0491_ ) );
NOR4_X1 \AXI4Interconnect/_1357_ ( .A1(\AXI4Interconnect/_0868_ ), .A2(\AXI4Interconnect/_0528_ ), .A3(\AXI4Interconnect/_0762_ ), .A4(fanout_net_4 ), .ZN(\AXI4Interconnect/_0492_ ) );
NOR4_X1 \AXI4Interconnect/_1358_ ( .A1(\AXI4Interconnect/_0868_ ), .A2(\AXI4Interconnect/_0528_ ), .A3(\AXI4Interconnect/_0763_ ), .A4(fanout_net_4 ), .ZN(\AXI4Interconnect/_0493_ ) );
BUF_X4 \AXI4Interconnect/_1359_ ( .A(\AXI4Interconnect/_0742_ ), .Z(\AXI4Interconnect/_0529_ ) );
NOR4_X1 \AXI4Interconnect/_1360_ ( .A1(\AXI4Interconnect/_0529_ ), .A2(\AXI4Interconnect/_0528_ ), .A3(\AXI4Interconnect/_0764_ ), .A4(fanout_net_4 ), .ZN(\AXI4Interconnect/_0494_ ) );
NOR4_X1 \AXI4Interconnect/_1361_ ( .A1(\AXI4Interconnect/_0529_ ), .A2(\AXI4Interconnect/_0528_ ), .A3(\AXI4Interconnect/_0765_ ), .A4(fanout_net_4 ), .ZN(\AXI4Interconnect/_0495_ ) );
NOR4_X1 \AXI4Interconnect/_1362_ ( .A1(\AXI4Interconnect/_0529_ ), .A2(\AXI4Interconnect/_0528_ ), .A3(\AXI4Interconnect/_0767_ ), .A4(fanout_net_4 ), .ZN(\AXI4Interconnect/_0496_ ) );
BUF_X4 \AXI4Interconnect/_1363_ ( .A(\AXI4Interconnect/_0622_ ), .Z(\AXI4Interconnect/_0530_ ) );
NOR4_X1 \AXI4Interconnect/_1364_ ( .A1(\AXI4Interconnect/_0529_ ), .A2(\AXI4Interconnect/_0530_ ), .A3(\AXI4Interconnect/_0768_ ), .A4(fanout_net_4 ), .ZN(\AXI4Interconnect/_0497_ ) );
NOR4_X1 \AXI4Interconnect/_1365_ ( .A1(\AXI4Interconnect/_0529_ ), .A2(\AXI4Interconnect/_0530_ ), .A3(\AXI4Interconnect/_0771_ ), .A4(fanout_net_4 ), .ZN(\AXI4Interconnect/_0498_ ) );
NOR4_X1 \AXI4Interconnect/_1366_ ( .A1(\AXI4Interconnect/_0529_ ), .A2(\AXI4Interconnect/_0530_ ), .A3(\AXI4Interconnect/_0772_ ), .A4(fanout_net_4 ), .ZN(\AXI4Interconnect/_0499_ ) );
NOR4_X1 \AXI4Interconnect/_1367_ ( .A1(\AXI4Interconnect/_0529_ ), .A2(\AXI4Interconnect/_0530_ ), .A3(\AXI4Interconnect/_0773_ ), .A4(fanout_net_4 ), .ZN(\AXI4Interconnect/_0501_ ) );
NOR4_X1 \AXI4Interconnect/_1368_ ( .A1(\AXI4Interconnect/_0529_ ), .A2(\AXI4Interconnect/_0530_ ), .A3(\AXI4Interconnect/_0774_ ), .A4(fanout_net_4 ), .ZN(\AXI4Interconnect/_0502_ ) );
NOR4_X1 \AXI4Interconnect/_1369_ ( .A1(\AXI4Interconnect/_0529_ ), .A2(\AXI4Interconnect/_0530_ ), .A3(\AXI4Interconnect/_0775_ ), .A4(fanout_net_4 ), .ZN(\AXI4Interconnect/_0503_ ) );
NOR4_X1 \AXI4Interconnect/_1370_ ( .A1(\AXI4Interconnect/_0529_ ), .A2(\AXI4Interconnect/_0530_ ), .A3(\AXI4Interconnect/_0776_ ), .A4(fanout_net_4 ), .ZN(\AXI4Interconnect/_0504_ ) );
BUF_X4 \AXI4Interconnect/_1371_ ( .A(\AXI4Interconnect/_0742_ ), .Z(\AXI4Interconnect/_0531_ ) );
NOR4_X1 \AXI4Interconnect/_1372_ ( .A1(\AXI4Interconnect/_0531_ ), .A2(\AXI4Interconnect/_0530_ ), .A3(\AXI4Interconnect/_0777_ ), .A4(fanout_net_4 ), .ZN(\AXI4Interconnect/_0505_ ) );
NOR4_X1 \AXI4Interconnect/_1373_ ( .A1(\AXI4Interconnect/_0531_ ), .A2(\AXI4Interconnect/_0530_ ), .A3(\AXI4Interconnect/_0778_ ), .A4(fanout_net_4 ), .ZN(\AXI4Interconnect/_0506_ ) );
NOR4_X1 \AXI4Interconnect/_1374_ ( .A1(\AXI4Interconnect/_0531_ ), .A2(\AXI4Interconnect/_0530_ ), .A3(\AXI4Interconnect/_0780_ ), .A4(fanout_net_4 ), .ZN(\AXI4Interconnect/_0507_ ) );
NOR4_X1 \AXI4Interconnect/_1375_ ( .A1(\AXI4Interconnect/_0531_ ), .A2(\AXI4Interconnect/_0618_ ), .A3(\AXI4Interconnect/_0781_ ), .A4(\AXI4Interconnect/_0004_ ), .ZN(\AXI4Interconnect/_0508_ ) );
NOR4_X1 \AXI4Interconnect/_1376_ ( .A1(\AXI4Interconnect/_0531_ ), .A2(\AXI4Interconnect/_0618_ ), .A3(\AXI4Interconnect/_0783_ ), .A4(\AXI4Interconnect/_0004_ ), .ZN(\AXI4Interconnect/_0509_ ) );
NOR4_X1 \AXI4Interconnect/_1377_ ( .A1(\AXI4Interconnect/_0531_ ), .A2(\AXI4Interconnect/_0618_ ), .A3(\AXI4Interconnect/_0784_ ), .A4(\AXI4Interconnect/_0004_ ), .ZN(\AXI4Interconnect/_0510_ ) );
NOR4_X1 \AXI4Interconnect/_1378_ ( .A1(\AXI4Interconnect/_0531_ ), .A2(\AXI4Interconnect/_0618_ ), .A3(\AXI4Interconnect/_0785_ ), .A4(\AXI4Interconnect/_0004_ ), .ZN(\AXI4Interconnect/_0512_ ) );
NOR4_X1 \AXI4Interconnect/_1379_ ( .A1(\AXI4Interconnect/_0531_ ), .A2(\AXI4Interconnect/_0618_ ), .A3(\AXI4Interconnect/_0786_ ), .A4(\AXI4Interconnect/_0004_ ), .ZN(\AXI4Interconnect/_0513_ ) );
INV_X1 \AXI4Interconnect/_1380_ ( .A(\AXI4Interconnect/_0611_ ), .ZN(\AXI4Interconnect/_0532_ ) );
CLKBUF_X2 \AXI4Interconnect/_1381_ ( .A(\AXI4Interconnect/_0532_ ), .Z(\AXI4Interconnect/_0533_ ) );
AND4_X1 \AXI4Interconnect/_1382_ ( .A1(\AXI4Interconnect/_0869_ ), .A2(\AXI4Interconnect/_0533_ ), .A3(\AXI4Interconnect/_0860_ ), .A4(\AXI4Interconnect/_0228_ ), .ZN(\AXI4Interconnect/_0523_ ) );
AND4_X1 \AXI4Interconnect/_1383_ ( .A1(\AXI4Interconnect/_0869_ ), .A2(\AXI4Interconnect/_0533_ ), .A3(\AXI4Interconnect/_0860_ ), .A4(\AXI4Interconnect/_0229_ ), .ZN(\AXI4Interconnect/_0524_ ) );
AND4_X1 \AXI4Interconnect/_1384_ ( .A1(\AXI4Interconnect/_0869_ ), .A2(\AXI4Interconnect/_0533_ ), .A3(\AXI4Interconnect/_0860_ ), .A4(\AXI4Interconnect/_0230_ ), .ZN(\AXI4Interconnect/_0525_ ) );
AND4_X1 \AXI4Interconnect/_1385_ ( .A1(\AXI4Interconnect/_0869_ ), .A2(\AXI4Interconnect/_0533_ ), .A3(\AXI4Interconnect/_0860_ ), .A4(\AXI4Interconnect/_0231_ ), .ZN(\AXI4Interconnect/_0526_ ) );
INV_X2 \AXI4Interconnect/_1386_ ( .A(\AXI4Interconnect/_0002_ ), .ZN(\AXI4Interconnect/_0534_ ) );
BUF_X4 \AXI4Interconnect/_1387_ ( .A(\AXI4Interconnect/_0534_ ), .Z(\AXI4Interconnect/_0535_ ) );
NOR2_X1 \AXI4Interconnect/_1388_ ( .A1(\AXI4Interconnect/_0535_ ), .A2(\AXI4Interconnect/_0792_ ), .ZN(\AXI4Interconnect/_0375_ ) );
NOR2_X1 \AXI4Interconnect/_1389_ ( .A1(\AXI4Interconnect/_0535_ ), .A2(\AXI4Interconnect/_0794_ ), .ZN(\AXI4Interconnect/_0386_ ) );
NOR2_X1 \AXI4Interconnect/_1390_ ( .A1(\AXI4Interconnect/_0535_ ), .A2(\AXI4Interconnect/_0796_ ), .ZN(\AXI4Interconnect/_0397_ ) );
NOR2_X1 \AXI4Interconnect/_1391_ ( .A1(\AXI4Interconnect/_0535_ ), .A2(\AXI4Interconnect/_0798_ ), .ZN(\AXI4Interconnect/_0400_ ) );
NOR2_X1 \AXI4Interconnect/_1392_ ( .A1(\AXI4Interconnect/_0535_ ), .A2(\AXI4Interconnect/_0800_ ), .ZN(\AXI4Interconnect/_0401_ ) );
NOR2_X1 \AXI4Interconnect/_1393_ ( .A1(\AXI4Interconnect/_0535_ ), .A2(\AXI4Interconnect/_0802_ ), .ZN(\AXI4Interconnect/_0402_ ) );
NOR2_X1 \AXI4Interconnect/_1394_ ( .A1(\AXI4Interconnect/_0535_ ), .A2(\AXI4Interconnect/_0804_ ), .ZN(\AXI4Interconnect/_0403_ ) );
BUF_X4 \AXI4Interconnect/_1395_ ( .A(\AXI4Interconnect/_0534_ ), .Z(\AXI4Interconnect/_0536_ ) );
NOR2_X1 \AXI4Interconnect/_1396_ ( .A1(\AXI4Interconnect/_0806_ ), .A2(\AXI4Interconnect/_0536_ ), .ZN(\AXI4Interconnect/_0404_ ) );
NOR2_X1 \AXI4Interconnect/_1397_ ( .A1(\AXI4Interconnect/_0809_ ), .A2(\AXI4Interconnect/_0536_ ), .ZN(\AXI4Interconnect/_0405_ ) );
NOR2_X1 \AXI4Interconnect/_1398_ ( .A1(\AXI4Interconnect/_0811_ ), .A2(\AXI4Interconnect/_0536_ ), .ZN(\AXI4Interconnect/_0406_ ) );
NOR2_X1 \AXI4Interconnect/_1399_ ( .A1(\AXI4Interconnect/_0535_ ), .A2(\AXI4Interconnect/_0813_ ), .ZN(\AXI4Interconnect/_0376_ ) );
NOR2_X1 \AXI4Interconnect/_1400_ ( .A1(\AXI4Interconnect/_0535_ ), .A2(\AXI4Interconnect/_0815_ ), .ZN(\AXI4Interconnect/_0377_ ) );
NOR2_X1 \AXI4Interconnect/_1401_ ( .A1(\AXI4Interconnect/_0817_ ), .A2(\AXI4Interconnect/_0536_ ), .ZN(\AXI4Interconnect/_0378_ ) );
NOR2_X1 \AXI4Interconnect/_1402_ ( .A1(\AXI4Interconnect/_0819_ ), .A2(\AXI4Interconnect/_0536_ ), .ZN(\AXI4Interconnect/_0379_ ) );
NOR2_X1 \AXI4Interconnect/_1403_ ( .A1(\AXI4Interconnect/_0535_ ), .A2(\AXI4Interconnect/_0821_ ), .ZN(\AXI4Interconnect/_0380_ ) );
BUF_X4 \AXI4Interconnect/_1404_ ( .A(\AXI4Interconnect/_0534_ ), .Z(\AXI4Interconnect/_0537_ ) );
NOR2_X1 \AXI4Interconnect/_1405_ ( .A1(\AXI4Interconnect/_0537_ ), .A2(\AXI4Interconnect/_0824_ ), .ZN(\AXI4Interconnect/_0381_ ) );
NOR2_X1 \AXI4Interconnect/_1406_ ( .A1(\AXI4Interconnect/_0537_ ), .A2(\AXI4Interconnect/_0826_ ), .ZN(\AXI4Interconnect/_0382_ ) );
NOR2_X1 \AXI4Interconnect/_1407_ ( .A1(\AXI4Interconnect/_0537_ ), .A2(\AXI4Interconnect/_0828_ ), .ZN(\AXI4Interconnect/_0383_ ) );
NOR2_X1 \AXI4Interconnect/_1408_ ( .A1(\AXI4Interconnect/_0537_ ), .A2(\AXI4Interconnect/_0830_ ), .ZN(\AXI4Interconnect/_0384_ ) );
NOR2_X1 \AXI4Interconnect/_1409_ ( .A1(\AXI4Interconnect/_0832_ ), .A2(\AXI4Interconnect/_0536_ ), .ZN(\AXI4Interconnect/_0385_ ) );
NOR2_X1 \AXI4Interconnect/_1410_ ( .A1(\AXI4Interconnect/_0537_ ), .A2(\AXI4Interconnect/_0834_ ), .ZN(\AXI4Interconnect/_0387_ ) );
NOR2_X1 \AXI4Interconnect/_1411_ ( .A1(\AXI4Interconnect/_0836_ ), .A2(\AXI4Interconnect/_0536_ ), .ZN(\AXI4Interconnect/_0388_ ) );
NOR2_X1 \AXI4Interconnect/_1412_ ( .A1(\AXI4Interconnect/_0838_ ), .A2(\AXI4Interconnect/_0534_ ), .ZN(\AXI4Interconnect/_0389_ ) );
NOR2_X1 \AXI4Interconnect/_1413_ ( .A1(\AXI4Interconnect/_0840_ ), .A2(\AXI4Interconnect/_0534_ ), .ZN(\AXI4Interconnect/_0390_ ) );
NOR2_X1 \AXI4Interconnect/_1414_ ( .A1(\AXI4Interconnect/_0842_ ), .A2(\AXI4Interconnect/_0534_ ), .ZN(\AXI4Interconnect/_0391_ ) );
NOR2_X1 \AXI4Interconnect/_1415_ ( .A1(\AXI4Interconnect/_0537_ ), .A2(\AXI4Interconnect/_0845_ ), .ZN(\AXI4Interconnect/_0392_ ) );
NOR2_X1 \AXI4Interconnect/_1416_ ( .A1(\AXI4Interconnect/_0537_ ), .A2(\AXI4Interconnect/_0848_ ), .ZN(\AXI4Interconnect/_0393_ ) );
NOR2_X1 \AXI4Interconnect/_1417_ ( .A1(\AXI4Interconnect/_0537_ ), .A2(\AXI4Interconnect/_0851_ ), .ZN(\AXI4Interconnect/_0394_ ) );
NOR2_X1 \AXI4Interconnect/_1418_ ( .A1(\AXI4Interconnect/_0537_ ), .A2(\AXI4Interconnect/_0853_ ), .ZN(\AXI4Interconnect/_0395_ ) );
NOR2_X1 \AXI4Interconnect/_1419_ ( .A1(\AXI4Interconnect/_0537_ ), .A2(\AXI4Interconnect/_0855_ ), .ZN(\AXI4Interconnect/_0396_ ) );
NOR2_X1 \AXI4Interconnect/_1420_ ( .A1(\AXI4Interconnect/_0536_ ), .A2(\AXI4Interconnect/_0857_ ), .ZN(\AXI4Interconnect/_0398_ ) );
NOR2_X1 \AXI4Interconnect/_1421_ ( .A1(\AXI4Interconnect/_0536_ ), .A2(\AXI4Interconnect/_0859_ ), .ZN(\AXI4Interconnect/_0399_ ) );
AND4_X1 \AXI4Interconnect/_1422_ ( .A1(\AXI4Interconnect/_0869_ ), .A2(\AXI4Interconnect/_0533_ ), .A3(\AXI4Interconnect/_0860_ ), .A4(\AXI4Interconnect/_0150_ ), .ZN(\AXI4Interconnect/_0445_ ) );
AND4_X1 \AXI4Interconnect/_1423_ ( .A1(\AXI4Interconnect/_0869_ ), .A2(\AXI4Interconnect/_0533_ ), .A3(\AXI4Interconnect/_0860_ ), .A4(\AXI4Interconnect/_0151_ ), .ZN(\AXI4Interconnect/_0446_ ) );
AND4_X1 \AXI4Interconnect/_1424_ ( .A1(\AXI4Interconnect/_0869_ ), .A2(\AXI4Interconnect/_0533_ ), .A3(\AXI4Interconnect/_0860_ ), .A4(\AXI4Interconnect/_0152_ ), .ZN(\AXI4Interconnect/_0447_ ) );
AND4_X1 \AXI4Interconnect/_1425_ ( .A1(\AXI4Interconnect/_0869_ ), .A2(\AXI4Interconnect/_0533_ ), .A3(\AXI4Interconnect/_0871_ ), .A4(\AXI4Interconnect/_0113_ ), .ZN(\AXI4Interconnect/_0408_ ) );
NOR2_X1 \AXI4Interconnect/_1426_ ( .A1(\AXI4Interconnect/_0779_ ), .A2(\AXI4Interconnect/_0114_ ), .ZN(\AXI4Interconnect/_0538_ ) );
NOR3_X1 \AXI4Interconnect/_1427_ ( .A1(\AXI4Interconnect/_0538_ ), .A2(\AXI4Interconnect/_0861_ ), .A3(\AXI4Interconnect/_0696_ ), .ZN(\AXI4Interconnect/_0409_ ) );
AND4_X1 \AXI4Interconnect/_1428_ ( .A1(\AXI4Interconnect/_0869_ ), .A2(\AXI4Interconnect/_0532_ ), .A3(\AXI4Interconnect/_0871_ ), .A4(\AXI4Interconnect/_0115_ ), .ZN(\AXI4Interconnect/_0410_ ) );
OR2_X1 \AXI4Interconnect/_1429_ ( .A1(\AXI4Interconnect/_0617_ ), .A2(\AXI4Interconnect/_0407_ ), .ZN(\AXI4Interconnect/_0539_ ) );
OAI21_X1 \AXI4Interconnect/_1430_ ( .A(\AXI4Interconnect/_0539_ ), .B1(\AXI4Interconnect/_0869_ ), .B2(\AXI4Interconnect/_0265_ ), .ZN(\AXI4Interconnect/_0540_ ) );
NOR2_X1 \AXI4Interconnect/_1431_ ( .A1(\AXI4Interconnect/_0540_ ), .A2(\AXI4Interconnect/_0614_ ), .ZN(\AXI4Interconnect/_0042_ ) );
NOR2_X2 \AXI4Interconnect/_1432_ ( .A1(\AXI4Interconnect/_0607_ ), .A2(\AXI4Interconnect/_0488_ ), .ZN(\AXI4Interconnect/_0541_ ) );
NOR2_X1 \AXI4Interconnect/_1433_ ( .A1(\AXI4Interconnect/_0869_ ), .A2(\AXI4Interconnect/_0340_ ), .ZN(\AXI4Interconnect/_0542_ ) );
NOR4_X1 \AXI4Interconnect/_1434_ ( .A1(\AXI4Interconnect/_0541_ ), .A2(\AXI4Interconnect/_0696_ ), .A3(\AXI4Interconnect/_0542_ ), .A4(\AXI4Interconnect/_0860_ ), .ZN(\AXI4Interconnect/_0079_ ) );
MUX2_X1 \AXI4Interconnect/_1435_ ( .A(\AXI4Interconnect/_0299_ ), .B(\AXI4Interconnect/_0444_ ), .S(\AXI4Interconnect/_0869_ ), .Z(\AXI4Interconnect/_0543_ ) );
AND2_X1 \AXI4Interconnect/_1436_ ( .A1(\AXI4Interconnect/_0543_ ), .A2(\AXI4Interconnect/_0690_ ), .ZN(\AXI4Interconnect/_0149_ ) );
MUX2_X1 \AXI4Interconnect/_1437_ ( .A(\AXI4Interconnect/_0373_ ), .B(\AXI4Interconnect/_0522_ ), .S(\AXI4Interconnect/_0869_ ), .Z(\AXI4Interconnect/_0544_ ) );
AND2_X1 \AXI4Interconnect/_1438_ ( .A1(\AXI4Interconnect/_0544_ ), .A2(\AXI4Interconnect/_0690_ ), .ZN(\AXI4Interconnect/_0227_ ) );
MUX2_X1 \AXI4Interconnect/_1439_ ( .A(\AXI4Interconnect/_0304_ ), .B(\AXI4Interconnect/_0452_ ), .S(\AXI4Interconnect/_0869_ ), .Z(\AXI4Interconnect/_0545_ ) );
AND2_X1 \AXI4Interconnect/_1440_ ( .A1(\AXI4Interconnect/_0545_ ), .A2(\AXI4Interconnect/_0690_ ), .ZN(\AXI4Interconnect/_0157_ ) );
NOR2_X1 \AXI4Interconnect/_1441_ ( .A1(\AXI4Interconnect/_0540_ ), .A2(\AXI4Interconnect/_0692_ ), .ZN(\AXI4Interconnect/_0112_ ) );
NOR4_X1 \AXI4Interconnect/_1442_ ( .A1(\AXI4Interconnect/_0541_ ), .A2(\AXI4Interconnect/_0696_ ), .A3(\AXI4Interconnect/_0542_ ), .A4(\AXI4Interconnect/_0779_ ), .ZN(\AXI4Interconnect/_0193_ ) );
INV_X32 \AXI4Interconnect/_1443_ ( .A(\AXI4Interconnect/_0153_ ), .ZN(\AXI4Interconnect/_0546_ ) );
NOR4_X1 \AXI4Interconnect/_1444_ ( .A1(\AXI4Interconnect/_0531_ ), .A2(\AXI4Interconnect/_0779_ ), .A3(\AXI4Interconnect/_0702_ ), .A4(\AXI4Interconnect/_0546_ ), .ZN(\AXI4Interconnect/_0300_ ) );
INV_X1 \AXI4Interconnect/_1445_ ( .A(\AXI4Interconnect/_0232_ ), .ZN(\AXI4Interconnect/_0547_ ) );
NOR4_X1 \AXI4Interconnect/_1446_ ( .A1(\AXI4Interconnect/_0531_ ), .A2(\AXI4Interconnect/_0779_ ), .A3(\AXI4Interconnect/_0702_ ), .A4(\AXI4Interconnect/_0547_ ), .ZN(\AXI4Interconnect/_0374_ ) );
INV_X1 \AXI4Interconnect/_1447_ ( .A(\AXI4Interconnect/_0154_ ), .ZN(\AXI4Interconnect/_0548_ ) );
OAI221_X1 \AXI4Interconnect/_1448_ ( .A(\AXI4Interconnect/_0005_ ), .B1(\AXI4Interconnect/_0873_ ), .B2(\AXI4Interconnect/_0872_ ), .C1(\AXI4Interconnect/_0700_ ), .C2(\AXI4Interconnect/_0548_ ), .ZN(\AXI4Interconnect/_0301_ ) );
INV_X32 \AXI4Interconnect/_1449_ ( .A(\AXI4Interconnect/_0043_ ), .ZN(\AXI4Interconnect/_0549_ ) );
INV_X32 \AXI4Interconnect/_1450_ ( .A(\AXI4Interconnect/_0116_ ), .ZN(\AXI4Interconnect/_0550_ ) );
MUX2_X1 \AXI4Interconnect/_1451_ ( .A(\AXI4Interconnect/_0549_ ), .B(\AXI4Interconnect/_0550_ ), .S(\AXI4Interconnect/_0871_ ), .Z(\AXI4Interconnect/_0551_ ) );
NOR2_X1 \AXI4Interconnect/_1452_ ( .A1(\AXI4Interconnect/_0807_ ), .A2(\AXI4Interconnect/_0551_ ), .ZN(\AXI4Interconnect/_0266_ ) );
NAND2_X4 \AXI4Interconnect/_1453_ ( .A1(\AXI4Interconnect/_0698_ ), .A2(\AXI4Interconnect/_0076_ ), .ZN(\AXI4Interconnect/_0552_ ) );
NAND2_X1 \AXI4Interconnect/_1454_ ( .A1(\AXI4Interconnect/_0871_ ), .A2(\AXI4Interconnect/_0190_ ), .ZN(\AXI4Interconnect/_0553_ ) );
NAND4_X1 \AXI4Interconnect/_1455_ ( .A1(\AXI4Interconnect/_0533_ ), .A2(\AXI4Interconnect/_0005_ ), .A3(\AXI4Interconnect/_0552_ ), .A4(\AXI4Interconnect/_0553_ ), .ZN(\AXI4Interconnect/_0337_ ) );
NOR4_X1 \AXI4Interconnect/_1456_ ( .A1(\AXI4Interconnect/_0696_ ), .A2(\AXI4Interconnect/_0618_ ), .A3(\AXI4Interconnect/_0546_ ), .A4(\AXI4Interconnect/_0004_ ), .ZN(\AXI4Interconnect/_0448_ ) );
NOR4_X1 \AXI4Interconnect/_1457_ ( .A1(\AXI4Interconnect/_0696_ ), .A2(\AXI4Interconnect/_0618_ ), .A3(\AXI4Interconnect/_0547_ ), .A4(\AXI4Interconnect/_0004_ ), .ZN(\AXI4Interconnect/_0527_ ) );
OAI221_X1 \AXI4Interconnect/_1458_ ( .A(\AXI4Interconnect/_0869_ ), .B1(\AXI4Interconnect/_0873_ ), .B2(\AXI4Interconnect/_0872_ ), .C1(\AXI4Interconnect/_0700_ ), .C2(\AXI4Interconnect/_0548_ ), .ZN(\AXI4Interconnect/_0449_ ) );
NOR2_X1 \AXI4Interconnect/_1459_ ( .A1(\AXI4Interconnect/_0536_ ), .A2(\AXI4Interconnect/_0551_ ), .ZN(\AXI4Interconnect/_0411_ ) );
NAND4_X1 \AXI4Interconnect/_1460_ ( .A1(\AXI4Interconnect/_0533_ ), .A2(\AXI4Interconnect/_0869_ ), .A3(\AXI4Interconnect/_0552_ ), .A4(\AXI4Interconnect/_0553_ ), .ZN(\AXI4Interconnect/_0485_ ) );
AND4_X1 \AXI4Interconnect/_1461_ ( .A1(\AXI4Interconnect/_0869_ ), .A2(\AXI4Interconnect/_0532_ ), .A3(\AXI4Interconnect/_0860_ ), .A4(\AXI4Interconnect/_0226_ ), .ZN(\AXI4Interconnect/_0521_ ) );
AOI211_X2 \AXI4Interconnect/_1462_ ( .A(\AXI4Interconnect/_0542_ ), .B(\AXI4Interconnect/_0541_ ), .C1(\AXI4Interconnect/_0552_ ), .C2(\AXI4Interconnect/_0553_ ), .ZN(\AXI4Interconnect/_0554_ ) );
AND2_X1 \AXI4Interconnect/_1463_ ( .A1(\AXI4Interconnect/_0873_ ), .A2(\AXI4Interconnect/_0872_ ), .ZN(\AXI4Interconnect/_0555_ ) );
INV_X1 \AXI4Interconnect/_1464_ ( .A(\AXI4Interconnect/_0555_ ), .ZN(\AXI4Interconnect/_0556_ ) );
NOR2_X1 \AXI4Interconnect/_1465_ ( .A1(\AXI4Interconnect/_0554_ ), .A2(\AXI4Interconnect/_0556_ ), .ZN(\AXI4Interconnect/_0557_ ) );
NOR2_X4 \AXI4Interconnect/_1466_ ( .A1(\AXI4Interconnect/_0043_ ), .A2(\AXI4Interconnect/_0116_ ), .ZN(\AXI4Interconnect/_0558_ ) );
INV_X2 \AXI4Interconnect/_1467_ ( .A(\AXI4Interconnect/_0558_ ), .ZN(\AXI4Interconnect/_0559_ ) );
OAI21_X1 \AXI4Interconnect/_1468_ ( .A(\AXI4Interconnect/_0611_ ), .B1(\AXI4Interconnect/_0559_ ), .B2(\AXI4Interconnect/_0153_ ), .ZN(\AXI4Interconnect/_0560_ ) );
NOR2_X4 \AXI4Interconnect/_1469_ ( .A1(\AXI4Interconnect/_0546_ ), .A2(\AXI4Interconnect/_0043_ ), .ZN(\AXI4Interconnect/_0561_ ) );
AOI21_X1 \AXI4Interconnect/_1470_ ( .A(\AXI4Interconnect/_0560_ ), .B1(\AXI4Interconnect/_0232_ ), .B2(\AXI4Interconnect/_0561_ ), .ZN(\AXI4Interconnect/_0562_ ) );
NOR2_X1 \AXI4Interconnect/_1471_ ( .A1(\AXI4Interconnect/_0557_ ), .A2(\AXI4Interconnect/_0562_ ), .ZN(\AXI4Interconnect/_0563_ ) );
AND3_X2 \AXI4Interconnect/_1472_ ( .A1(\AXI4Interconnect/_0544_ ), .A2(\AXI4Interconnect/_0232_ ), .A3(\AXI4Interconnect/_0690_ ), .ZN(\AXI4Interconnect/_0564_ ) );
INV_X1 \AXI4Interconnect/_1473_ ( .A(\AXI4Interconnect/_0872_ ), .ZN(\AXI4Interconnect/_0565_ ) );
OR3_X1 \AXI4Interconnect/_1474_ ( .A1(\AXI4Interconnect/_0564_ ), .A2(\AXI4Interconnect/_0873_ ), .A3(\AXI4Interconnect/_0565_ ), .ZN(\AXI4Interconnect/_0566_ ) );
AOI21_X1 \AXI4Interconnect/_1475_ ( .A(\AXI4Interconnect/_0870_ ), .B1(\AXI4Interconnect/_0563_ ), .B2(\AXI4Interconnect/_0566_ ), .ZN(\AXI4Interconnect/_0006_ ) );
INV_X1 \AXI4Interconnect/_1476_ ( .A(\AXI4Interconnect/_0564_ ), .ZN(\AXI4Interconnect/_0567_ ) );
NOR3_X1 \AXI4Interconnect/_1477_ ( .A1(\AXI4Interconnect/_0567_ ), .A2(\AXI4Interconnect/_0873_ ), .A3(\AXI4Interconnect/_0565_ ), .ZN(\AXI4Interconnect/_0568_ ) );
NAND3_X1 \AXI4Interconnect/_1478_ ( .A1(\AXI4Interconnect/_0545_ ), .A2(\AXI4Interconnect/_0154_ ), .A3(\AXI4Interconnect/_0690_ ), .ZN(\AXI4Interconnect/_0569_ ) );
AND3_X1 \AXI4Interconnect/_1479_ ( .A1(\AXI4Interconnect/_0569_ ), .A2(\AXI4Interconnect/_0873_ ), .A3(\AXI4Interconnect/_0565_ ), .ZN(\AXI4Interconnect/_0570_ ) );
AOI21_X1 \AXI4Interconnect/_1480_ ( .A(\AXI4Interconnect/_0560_ ), .B1(\AXI4Interconnect/_0547_ ), .B2(\AXI4Interconnect/_0561_ ), .ZN(\AXI4Interconnect/_0571_ ) );
NOR4_X1 \AXI4Interconnect/_1481_ ( .A1(\AXI4Interconnect/_0568_ ), .A2(\AXI4Interconnect/_0557_ ), .A3(\AXI4Interconnect/_0570_ ), .A4(\AXI4Interconnect/_0571_ ), .ZN(\AXI4Interconnect/_0572_ ) );
NOR2_X1 \AXI4Interconnect/_1482_ ( .A1(\AXI4Interconnect/_0572_ ), .A2(\AXI4Interconnect/_0870_ ), .ZN(\AXI4Interconnect/_0007_ ) );
NAND2_X1 \AXI4Interconnect/_1483_ ( .A1(\AXI4Interconnect/_0696_ ), .A2(\AXI4Interconnect/_0549_ ), .ZN(\AXI4Interconnect/_0573_ ) );
AOI21_X1 \AXI4Interconnect/_1484_ ( .A(\AXI4Interconnect/_0870_ ), .B1(\AXI4Interconnect/_0692_ ), .B2(\AXI4Interconnect/_0573_ ), .ZN(\AXI4Interconnect/_0008_ ) );
AND2_X1 \AXI4Interconnect/_1485_ ( .A1(\AXI4Interconnect/_0561_ ), .A2(\AXI4Interconnect/_0610_ ), .ZN(\AXI4Interconnect/_0574_ ) );
NAND4_X1 \AXI4Interconnect/_1486_ ( .A1(\AXI4Interconnect/_0574_ ), .A2(\AXI4Interconnect/_0735_ ), .A3(\AXI4Interconnect/_0134_ ), .A4(\AXI4Interconnect/_0558_ ), .ZN(\AXI4Interconnect/_0575_ ) );
NOR3_X1 \AXI4Interconnect/_1487_ ( .A1(\AXI4Interconnect/_0843_ ), .A2(\AXI4Interconnect/_0549_ ), .A3(\AXI4Interconnect/_0026_ ), .ZN(\AXI4Interconnect/_0576_ ) );
NOR3_X2 \AXI4Interconnect/_1488_ ( .A1(\AXI4Interconnect/_0844_ ), .A2(\AXI4Interconnect/_0096_ ), .A3(\AXI4Interconnect/_0043_ ), .ZN(\AXI4Interconnect/_0577_ ) );
OAI211_X2 \AXI4Interconnect/_1489_ ( .A(\AXI4Interconnect/_0611_ ), .B(\AXI4Interconnect/_0559_ ), .C1(\AXI4Interconnect/_0576_ ), .C2(\AXI4Interconnect/_0577_ ), .ZN(\AXI4Interconnect/_0578_ ) );
NAND2_X1 \AXI4Interconnect/_1490_ ( .A1(\AXI4Interconnect/_0575_ ), .A2(\AXI4Interconnect/_0578_ ), .ZN(\AXI4Interconnect/_0579_ ) );
NAND3_X1 \AXI4Interconnect/_1491_ ( .A1(\AXI4Interconnect/_0847_ ), .A2(\AXI4Interconnect/_0850_ ), .A3(\AXI4Interconnect/_0549_ ), .ZN(\AXI4Interconnect/_0580_ ) );
AND3_X2 \AXI4Interconnect/_1492_ ( .A1(\AXI4Interconnect/_0580_ ), .A2(\AXI4Interconnect/_0559_ ), .A3(\AXI4Interconnect/_0611_ ), .ZN(\AXI4Interconnect/_0581_ ) );
NAND3_X1 \AXI4Interconnect/_1493_ ( .A1(\AXI4Interconnect/_0846_ ), .A2(\AXI4Interconnect/_0849_ ), .A3(\AXI4Interconnect/_0043_ ), .ZN(\AXI4Interconnect/_0582_ ) );
NAND2_X1 \AXI4Interconnect/_1494_ ( .A1(\AXI4Interconnect/_0581_ ), .A2(\AXI4Interconnect/_0582_ ), .ZN(\AXI4Interconnect/_0583_ ) );
NAND2_X1 \AXI4Interconnect/_1495_ ( .A1(\AXI4Interconnect/_0737_ ), .A2(\AXI4Interconnect/_0738_ ), .ZN(\AXI4Interconnect/_0584_ ) );
NAND3_X1 \AXI4Interconnect/_1496_ ( .A1(\AXI4Interconnect/_0574_ ), .A2(\AXI4Interconnect/_0558_ ), .A3(\AXI4Interconnect/_0584_ ), .ZN(\AXI4Interconnect/_0585_ ) );
AND3_X2 \AXI4Interconnect/_1497_ ( .A1(\AXI4Interconnect/_0579_ ), .A2(\AXI4Interconnect/_0583_ ), .A3(\AXI4Interconnect/_0585_ ), .ZN(\AXI4Interconnect/_0586_ ) );
NAND4_X1 \AXI4Interconnect/_1498_ ( .A1(\AXI4Interconnect/_0740_ ), .A2(\AXI4Interconnect/_0741_ ), .A3(\AXI4Interconnect/_0745_ ), .A4(\AXI4Interconnect/_0746_ ), .ZN(\AXI4Interconnect/_0587_ ) );
AOI21_X1 \AXI4Interconnect/_1499_ ( .A(\AXI4Interconnect/_0559_ ), .B1(\AXI4Interconnect/_0587_ ), .B2(\AXI4Interconnect/_0153_ ), .ZN(\AXI4Interconnect/_0588_ ) );
OR4_X4 \AXI4Interconnect/_1500_ ( .A1(\AXI4Interconnect/_0100_ ), .A2(\AXI4Interconnect/_0550_ ), .A3(\AXI4Interconnect/_0101_ ), .A4(\AXI4Interconnect/_0104_ ), .ZN(\AXI4Interconnect/_0589_ ) );
OR3_X4 \AXI4Interconnect/_1501_ ( .A1(\AXI4Interconnect/_0589_ ), .A2(\AXI4Interconnect/_0103_ ), .A3(\AXI4Interconnect/_0043_ ), .ZN(\AXI4Interconnect/_0590_ ) );
OR4_X1 \AXI4Interconnect/_1502_ ( .A1(\AXI4Interconnect/_0030_ ), .A2(\AXI4Interconnect/_0549_ ), .A3(\AXI4Interconnect/_0031_ ), .A4(\AXI4Interconnect/_0034_ ), .ZN(\AXI4Interconnect/_0591_ ) );
OAI21_X2 \AXI4Interconnect/_1503_ ( .A(\AXI4Interconnect/_0590_ ), .B1(\AXI4Interconnect/_0033_ ), .B2(\AXI4Interconnect/_0591_ ), .ZN(\AXI4Interconnect/_0592_ ) );
OAI21_X1 \AXI4Interconnect/_1504_ ( .A(\AXI4Interconnect/_0586_ ), .B1(\AXI4Interconnect/_0588_ ), .B2(\AXI4Interconnect/_0592_ ), .ZN(\AXI4Interconnect/_0593_ ) );
NOR4_X1 \AXI4Interconnect/_1505_ ( .A1(\AXI4Interconnect/_0092_ ), .A2(\AXI4Interconnect/_0093_ ), .A3(\AXI4Interconnect/_0094_ ), .A4(\AXI4Interconnect/_0095_ ), .ZN(\AXI4Interconnect/_0594_ ) );
NOR4_X4 \AXI4Interconnect/_1506_ ( .A1(\AXI4Interconnect/_0087_ ), .A2(\AXI4Interconnect/_0088_ ), .A3(\AXI4Interconnect/_0089_ ), .A4(\AXI4Interconnect/_0090_ ), .ZN(\AXI4Interconnect/_0595_ ) );
AND4_X1 \AXI4Interconnect/_1507_ ( .A1(\AXI4Interconnect/_0549_ ), .A2(\AXI4Interconnect/_0594_ ), .A3(\AXI4Interconnect/_0595_ ), .A4(\AXI4Interconnect/_0116_ ), .ZN(\AXI4Interconnect/_0596_ ) );
NOR4_X4 \AXI4Interconnect/_1508_ ( .A1(\AXI4Interconnect/_0129_ ), .A2(\AXI4Interconnect/_0130_ ), .A3(\AXI4Interconnect/_0131_ ), .A4(\AXI4Interconnect/_0132_ ), .ZN(\AXI4Interconnect/_0597_ ) );
NOR4_X4 \AXI4Interconnect/_1509_ ( .A1(\AXI4Interconnect/_0124_ ), .A2(\AXI4Interconnect/_0125_ ), .A3(\AXI4Interconnect/_0126_ ), .A4(\AXI4Interconnect/_0127_ ), .ZN(\AXI4Interconnect/_0598_ ) );
NAND2_X1 \AXI4Interconnect/_1510_ ( .A1(\AXI4Interconnect/_0597_ ), .A2(\AXI4Interconnect/_0598_ ), .ZN(\AXI4Interconnect/_0599_ ) );
AOI21_X1 \AXI4Interconnect/_1511_ ( .A(\AXI4Interconnect/_0559_ ), .B1(\AXI4Interconnect/_0599_ ), .B2(\AXI4Interconnect/_0153_ ), .ZN(\AXI4Interconnect/_0600_ ) );
NOR3_X1 \AXI4Interconnect/_1512_ ( .A1(\AXI4Interconnect/_0549_ ), .A2(\AXI4Interconnect/_0024_ ), .A3(\AXI4Interconnect/_0025_ ), .ZN(\AXI4Interconnect/_0601_ ) );
OR4_X4 \AXI4Interconnect/_1513_ ( .A1(\AXI4Interconnect/_0019_ ), .A2(\AXI4Interconnect/_0020_ ), .A3(\AXI4Interconnect/_0022_ ), .A4(\AXI4Interconnect/_0023_ ), .ZN(\AXI4Interconnect/_0602_ ) );
NOR3_X1 \AXI4Interconnect/_1514_ ( .A1(\AXI4Interconnect/_0602_ ), .A2(\AXI4Interconnect/_0017_ ), .A3(\AXI4Interconnect/_0018_ ), .ZN(\AXI4Interconnect/_0603_ ) );
AOI211_X4 \AXI4Interconnect/_1515_ ( .A(\AXI4Interconnect/_0596_ ), .B(\AXI4Interconnect/_0600_ ), .C1(\AXI4Interconnect/_0601_ ), .C2(\AXI4Interconnect/_0603_ ), .ZN(\AXI4Interconnect/_0604_ ) );
OAI21_X1 \AXI4Interconnect/_1516_ ( .A(\AXI4Interconnect/_0696_ ), .B1(\AXI4Interconnect/_0593_ ), .B2(\AXI4Interconnect/_0604_ ), .ZN(\AXI4Interconnect/_0605_ ) );
AOI21_X1 \AXI4Interconnect/_1517_ ( .A(\AXI4Interconnect/_0870_ ), .B1(\AXI4Interconnect/_0605_ ), .B2(\AXI4Interconnect/_0534_ ), .ZN(\AXI4Interconnect/_0009_ ) );
DFF_X1 \AXI4Interconnect/_1518_ ( .D(\AXI4Interconnect/_0877_ ), .CK(clock ), .Q(\AXI4Interconnect/state [0] ), .QN(\AXI4Interconnect/_0875_ ) );
DFF_X1 \AXI4Interconnect/_1519_ ( .D(\AXI4Interconnect/_0878_ ), .CK(clock ), .Q(\AXI4Interconnect/state [1] ), .QN(\AXI4Interconnect/_0874_ ) );
DFF_X1 \AXI4Interconnect/_1520_ ( .D(\AXI4Interconnect/_0879_ ), .CK(clock ), .Q(\AXI4Interconnect/selectedReg ), .QN(\AXI4Interconnect/_0000_ ) );
DFF_X1 \AXI4Interconnect/_1521_ ( .D(\AXI4Interconnect/_0880_ ), .CK(clock ), .Q(\AXI4Interconnect/outSelect ), .QN(\AXI4Interconnect/_0001_ ) );
LOGIC0_X1 \AXI4Interconnect/_1522_ ( .Z(\AXI4Interconnect/_0876_ ) );
BUF_X1 \AXI4Interconnect/_1523_ ( .A(\AXI4Interconnect/_GEN_13 ), .Z(\io_master_arburst [0] ) );
BUF_X1 \AXI4Interconnect/_1524_ ( .A(\AXI4Interconnect/_0876_ ), .Z(\io_master_arburst [1] ) );
BUF_X1 \AXI4Interconnect/_1525_ ( .A(\AXI4Interconnect/_GEN_14 ), .Z(\io_master_awburst [0] ) );
BUF_X1 \AXI4Interconnect/_1526_ ( .A(\AXI4Interconnect/_0876_ ), .Z(\io_master_awburst [1] ) );
BUF_X1 \AXI4Interconnect/_1527_ ( .A(\AXI4Interconnect/state [1] ), .Z(\AXI4Interconnect/_0873_ ) );
BUF_X1 \AXI4Interconnect/_1528_ ( .A(\AXI4Interconnect/state [0] ), .Z(\AXI4Interconnect/_0872_ ) );
BUF_X1 \AXI4Interconnect/_1529_ ( .A(\_CLINT_io_rresp [0] ), .Z(\AXI4Interconnect/_0338_ ) );
BUF_X1 \AXI4Interconnect/_1530_ ( .A(\io_master_rresp [0] ), .Z(\AXI4Interconnect/_0486_ ) );
BUF_X1 \AXI4Interconnect/_1531_ ( .A(\AXI4Interconnect/outSelect ), .Z(\AXI4Interconnect/_0869_ ) );
BUF_X1 \AXI4Interconnect/_1532_ ( .A(\AXI4Interconnect/_0000_ ), .Z(\AXI4Interconnect/_0004_ ) );
BUF_X1 \AXI4Interconnect/_1533_ ( .A(\AXI4Interconnect/_0077_ ), .Z(\_AXI4Interconnect_io_fanIn_0_rresp [0] ) );
BUF_X1 \AXI4Interconnect/_1534_ ( .A(\_CLINT_io_rresp [1] ), .Z(\AXI4Interconnect/_0339_ ) );
BUF_X1 \AXI4Interconnect/_1535_ ( .A(\io_master_rresp [1] ), .Z(\AXI4Interconnect/_0487_ ) );
BUF_X1 \AXI4Interconnect/_1536_ ( .A(\AXI4Interconnect/_0078_ ), .Z(\_AXI4Interconnect_io_fanIn_0_rresp [1] ) );
BUF_X1 \AXI4Interconnect/_1537_ ( .A(\_CLINT_io_rdata [0] ), .Z(\AXI4Interconnect/_0305_ ) );
BUF_X1 \AXI4Interconnect/_1538_ ( .A(\io_master_rdata [0] ), .Z(\AXI4Interconnect/_0453_ ) );
BUF_X1 \AXI4Interconnect/_1539_ ( .A(\AXI4Interconnect/_0044_ ), .Z(\_AXI4Interconnect_io_fanIn_0_rdata [0] ) );
BUF_X1 \AXI4Interconnect/_1540_ ( .A(\_CLINT_io_rdata [1] ), .Z(\AXI4Interconnect/_0316_ ) );
BUF_X1 \AXI4Interconnect/_1541_ ( .A(\io_master_rdata [1] ), .Z(\AXI4Interconnect/_0464_ ) );
BUF_X1 \AXI4Interconnect/_1542_ ( .A(\AXI4Interconnect/_0055_ ), .Z(\_AXI4Interconnect_io_fanIn_0_rdata [1] ) );
BUF_X1 \AXI4Interconnect/_1543_ ( .A(\_CLINT_io_rdata [2] ), .Z(\AXI4Interconnect/_0327_ ) );
BUF_X1 \AXI4Interconnect/_1544_ ( .A(\io_master_rdata [2] ), .Z(\AXI4Interconnect/_0475_ ) );
BUF_X1 \AXI4Interconnect/_1545_ ( .A(\AXI4Interconnect/_0066_ ), .Z(\_AXI4Interconnect_io_fanIn_0_rdata [2] ) );
BUF_X1 \AXI4Interconnect/_1546_ ( .A(\_CLINT_io_rdata [3] ), .Z(\AXI4Interconnect/_0330_ ) );
BUF_X1 \AXI4Interconnect/_1547_ ( .A(\io_master_rdata [3] ), .Z(\AXI4Interconnect/_0478_ ) );
BUF_X1 \AXI4Interconnect/_1548_ ( .A(\AXI4Interconnect/_0069_ ), .Z(\_AXI4Interconnect_io_fanIn_0_rdata [3] ) );
BUF_X1 \AXI4Interconnect/_1549_ ( .A(\_CLINT_io_rdata [4] ), .Z(\AXI4Interconnect/_0331_ ) );
BUF_X1 \AXI4Interconnect/_1550_ ( .A(\io_master_rdata [4] ), .Z(\AXI4Interconnect/_0479_ ) );
BUF_X1 \AXI4Interconnect/_1551_ ( .A(\AXI4Interconnect/_0070_ ), .Z(\_AXI4Interconnect_io_fanIn_0_rdata [4] ) );
BUF_X1 \AXI4Interconnect/_1552_ ( .A(\_CLINT_io_rdata [5] ), .Z(\AXI4Interconnect/_0332_ ) );
BUF_X1 \AXI4Interconnect/_1553_ ( .A(\io_master_rdata [5] ), .Z(\AXI4Interconnect/_0480_ ) );
BUF_X1 \AXI4Interconnect/_1554_ ( .A(\AXI4Interconnect/_0071_ ), .Z(\_AXI4Interconnect_io_fanIn_0_rdata [5] ) );
BUF_X1 \AXI4Interconnect/_1555_ ( .A(\_CLINT_io_rdata [6] ), .Z(\AXI4Interconnect/_0333_ ) );
BUF_X1 \AXI4Interconnect/_1556_ ( .A(\io_master_rdata [6] ), .Z(\AXI4Interconnect/_0481_ ) );
BUF_X1 \AXI4Interconnect/_1557_ ( .A(\AXI4Interconnect/_0072_ ), .Z(\_AXI4Interconnect_io_fanIn_0_rdata [6] ) );
BUF_X1 \AXI4Interconnect/_1558_ ( .A(\_CLINT_io_rdata [7] ), .Z(\AXI4Interconnect/_0334_ ) );
BUF_X1 \AXI4Interconnect/_1559_ ( .A(\io_master_rdata [7] ), .Z(\AXI4Interconnect/_0482_ ) );
BUF_X1 \AXI4Interconnect/_1560_ ( .A(\AXI4Interconnect/_0073_ ), .Z(\_AXI4Interconnect_io_fanIn_0_rdata [7] ) );
BUF_X1 \AXI4Interconnect/_1561_ ( .A(\_CLINT_io_rdata [8] ), .Z(\AXI4Interconnect/_0335_ ) );
BUF_X1 \AXI4Interconnect/_1562_ ( .A(\io_master_rdata [8] ), .Z(\AXI4Interconnect/_0483_ ) );
BUF_X1 \AXI4Interconnect/_1563_ ( .A(\AXI4Interconnect/_0074_ ), .Z(\_AXI4Interconnect_io_fanIn_0_rdata [8] ) );
BUF_X1 \AXI4Interconnect/_1564_ ( .A(\_CLINT_io_rdata [9] ), .Z(\AXI4Interconnect/_0336_ ) );
BUF_X1 \AXI4Interconnect/_1565_ ( .A(\io_master_rdata [9] ), .Z(\AXI4Interconnect/_0484_ ) );
BUF_X1 \AXI4Interconnect/_1566_ ( .A(\AXI4Interconnect/_0075_ ), .Z(\_AXI4Interconnect_io_fanIn_0_rdata [9] ) );
BUF_X1 \AXI4Interconnect/_1567_ ( .A(\_CLINT_io_rdata [10] ), .Z(\AXI4Interconnect/_0306_ ) );
BUF_X1 \AXI4Interconnect/_1568_ ( .A(\io_master_rdata [10] ), .Z(\AXI4Interconnect/_0454_ ) );
BUF_X1 \AXI4Interconnect/_1569_ ( .A(\AXI4Interconnect/_0045_ ), .Z(\_AXI4Interconnect_io_fanIn_0_rdata [10] ) );
BUF_X1 \AXI4Interconnect/_1570_ ( .A(\_CLINT_io_rdata [11] ), .Z(\AXI4Interconnect/_0307_ ) );
BUF_X1 \AXI4Interconnect/_1571_ ( .A(\io_master_rdata [11] ), .Z(\AXI4Interconnect/_0455_ ) );
BUF_X1 \AXI4Interconnect/_1572_ ( .A(\AXI4Interconnect/_0046_ ), .Z(\_AXI4Interconnect_io_fanIn_0_rdata [11] ) );
BUF_X1 \AXI4Interconnect/_1573_ ( .A(\_CLINT_io_rdata [12] ), .Z(\AXI4Interconnect/_0308_ ) );
BUF_X1 \AXI4Interconnect/_1574_ ( .A(\io_master_rdata [12] ), .Z(\AXI4Interconnect/_0456_ ) );
BUF_X1 \AXI4Interconnect/_1575_ ( .A(\AXI4Interconnect/_0047_ ), .Z(\_AXI4Interconnect_io_fanIn_0_rdata [12] ) );
BUF_X1 \AXI4Interconnect/_1576_ ( .A(\_CLINT_io_rdata [13] ), .Z(\AXI4Interconnect/_0309_ ) );
BUF_X1 \AXI4Interconnect/_1577_ ( .A(\io_master_rdata [13] ), .Z(\AXI4Interconnect/_0457_ ) );
BUF_X1 \AXI4Interconnect/_1578_ ( .A(\AXI4Interconnect/_0048_ ), .Z(\_AXI4Interconnect_io_fanIn_0_rdata [13] ) );
BUF_X1 \AXI4Interconnect/_1579_ ( .A(\_CLINT_io_rdata [14] ), .Z(\AXI4Interconnect/_0310_ ) );
BUF_X1 \AXI4Interconnect/_1580_ ( .A(\io_master_rdata [14] ), .Z(\AXI4Interconnect/_0458_ ) );
BUF_X1 \AXI4Interconnect/_1581_ ( .A(\AXI4Interconnect/_0049_ ), .Z(\_AXI4Interconnect_io_fanIn_0_rdata [14] ) );
BUF_X1 \AXI4Interconnect/_1582_ ( .A(\_CLINT_io_rdata [15] ), .Z(\AXI4Interconnect/_0311_ ) );
BUF_X1 \AXI4Interconnect/_1583_ ( .A(\io_master_rdata [15] ), .Z(\AXI4Interconnect/_0459_ ) );
BUF_X1 \AXI4Interconnect/_1584_ ( .A(\AXI4Interconnect/_0050_ ), .Z(\_AXI4Interconnect_io_fanIn_0_rdata [15] ) );
BUF_X1 \AXI4Interconnect/_1585_ ( .A(\_CLINT_io_rdata [16] ), .Z(\AXI4Interconnect/_0312_ ) );
BUF_X1 \AXI4Interconnect/_1586_ ( .A(\io_master_rdata [16] ), .Z(\AXI4Interconnect/_0460_ ) );
BUF_X1 \AXI4Interconnect/_1587_ ( .A(\AXI4Interconnect/_0051_ ), .Z(\_AXI4Interconnect_io_fanIn_0_rdata [16] ) );
BUF_X1 \AXI4Interconnect/_1588_ ( .A(\_CLINT_io_rdata [17] ), .Z(\AXI4Interconnect/_0313_ ) );
BUF_X1 \AXI4Interconnect/_1589_ ( .A(\io_master_rdata [17] ), .Z(\AXI4Interconnect/_0461_ ) );
BUF_X1 \AXI4Interconnect/_1590_ ( .A(\AXI4Interconnect/_0052_ ), .Z(\_AXI4Interconnect_io_fanIn_0_rdata [17] ) );
BUF_X1 \AXI4Interconnect/_1591_ ( .A(\_CLINT_io_rdata [18] ), .Z(\AXI4Interconnect/_0314_ ) );
BUF_X1 \AXI4Interconnect/_1592_ ( .A(\io_master_rdata [18] ), .Z(\AXI4Interconnect/_0462_ ) );
BUF_X1 \AXI4Interconnect/_1593_ ( .A(\AXI4Interconnect/_0053_ ), .Z(\_AXI4Interconnect_io_fanIn_0_rdata [18] ) );
BUF_X1 \AXI4Interconnect/_1594_ ( .A(\_CLINT_io_rdata [19] ), .Z(\AXI4Interconnect/_0315_ ) );
BUF_X1 \AXI4Interconnect/_1595_ ( .A(\io_master_rdata [19] ), .Z(\AXI4Interconnect/_0463_ ) );
BUF_X1 \AXI4Interconnect/_1596_ ( .A(\AXI4Interconnect/_0054_ ), .Z(\_AXI4Interconnect_io_fanIn_0_rdata [19] ) );
BUF_X1 \AXI4Interconnect/_1597_ ( .A(\_CLINT_io_rdata [20] ), .Z(\AXI4Interconnect/_0317_ ) );
BUF_X1 \AXI4Interconnect/_1598_ ( .A(\io_master_rdata [20] ), .Z(\AXI4Interconnect/_0465_ ) );
BUF_X1 \AXI4Interconnect/_1599_ ( .A(\AXI4Interconnect/_0056_ ), .Z(\_AXI4Interconnect_io_fanIn_0_rdata [20] ) );
BUF_X1 \AXI4Interconnect/_1600_ ( .A(\_CLINT_io_rdata [21] ), .Z(\AXI4Interconnect/_0318_ ) );
BUF_X1 \AXI4Interconnect/_1601_ ( .A(\io_master_rdata [21] ), .Z(\AXI4Interconnect/_0466_ ) );
BUF_X1 \AXI4Interconnect/_1602_ ( .A(\AXI4Interconnect/_0057_ ), .Z(\_AXI4Interconnect_io_fanIn_0_rdata [21] ) );
BUF_X1 \AXI4Interconnect/_1603_ ( .A(\_CLINT_io_rdata [22] ), .Z(\AXI4Interconnect/_0319_ ) );
BUF_X1 \AXI4Interconnect/_1604_ ( .A(\io_master_rdata [22] ), .Z(\AXI4Interconnect/_0467_ ) );
BUF_X1 \AXI4Interconnect/_1605_ ( .A(\AXI4Interconnect/_0058_ ), .Z(\_AXI4Interconnect_io_fanIn_0_rdata [22] ) );
BUF_X1 \AXI4Interconnect/_1606_ ( .A(\_CLINT_io_rdata [23] ), .Z(\AXI4Interconnect/_0320_ ) );
BUF_X1 \AXI4Interconnect/_1607_ ( .A(\io_master_rdata [23] ), .Z(\AXI4Interconnect/_0468_ ) );
BUF_X1 \AXI4Interconnect/_1608_ ( .A(\AXI4Interconnect/_0059_ ), .Z(\_AXI4Interconnect_io_fanIn_0_rdata [23] ) );
BUF_X1 \AXI4Interconnect/_1609_ ( .A(\_CLINT_io_rdata [24] ), .Z(\AXI4Interconnect/_0321_ ) );
BUF_X1 \AXI4Interconnect/_1610_ ( .A(\io_master_rdata [24] ), .Z(\AXI4Interconnect/_0469_ ) );
BUF_X1 \AXI4Interconnect/_1611_ ( .A(\AXI4Interconnect/_0060_ ), .Z(\_AXI4Interconnect_io_fanIn_0_rdata [24] ) );
BUF_X1 \AXI4Interconnect/_1612_ ( .A(\_CLINT_io_rdata [25] ), .Z(\AXI4Interconnect/_0322_ ) );
BUF_X1 \AXI4Interconnect/_1613_ ( .A(\io_master_rdata [25] ), .Z(\AXI4Interconnect/_0470_ ) );
BUF_X1 \AXI4Interconnect/_1614_ ( .A(\AXI4Interconnect/_0061_ ), .Z(\_AXI4Interconnect_io_fanIn_0_rdata [25] ) );
BUF_X1 \AXI4Interconnect/_1615_ ( .A(\_CLINT_io_rdata [26] ), .Z(\AXI4Interconnect/_0323_ ) );
BUF_X1 \AXI4Interconnect/_1616_ ( .A(\io_master_rdata [26] ), .Z(\AXI4Interconnect/_0471_ ) );
BUF_X1 \AXI4Interconnect/_1617_ ( .A(\AXI4Interconnect/_0062_ ), .Z(\_AXI4Interconnect_io_fanIn_0_rdata [26] ) );
BUF_X1 \AXI4Interconnect/_1618_ ( .A(\_CLINT_io_rdata [27] ), .Z(\AXI4Interconnect/_0324_ ) );
BUF_X1 \AXI4Interconnect/_1619_ ( .A(\io_master_rdata [27] ), .Z(\AXI4Interconnect/_0472_ ) );
BUF_X1 \AXI4Interconnect/_1620_ ( .A(\AXI4Interconnect/_0063_ ), .Z(\_AXI4Interconnect_io_fanIn_0_rdata [27] ) );
BUF_X1 \AXI4Interconnect/_1621_ ( .A(\_CLINT_io_rdata [28] ), .Z(\AXI4Interconnect/_0325_ ) );
BUF_X1 \AXI4Interconnect/_1622_ ( .A(\io_master_rdata [28] ), .Z(\AXI4Interconnect/_0473_ ) );
BUF_X1 \AXI4Interconnect/_1623_ ( .A(\AXI4Interconnect/_0064_ ), .Z(\_AXI4Interconnect_io_fanIn_0_rdata [28] ) );
BUF_X1 \AXI4Interconnect/_1624_ ( .A(\_CLINT_io_rdata [29] ), .Z(\AXI4Interconnect/_0326_ ) );
BUF_X1 \AXI4Interconnect/_1625_ ( .A(\io_master_rdata [29] ), .Z(\AXI4Interconnect/_0474_ ) );
BUF_X1 \AXI4Interconnect/_1626_ ( .A(\AXI4Interconnect/_0065_ ), .Z(\_AXI4Interconnect_io_fanIn_0_rdata [29] ) );
BUF_X1 \AXI4Interconnect/_1627_ ( .A(\_CLINT_io_rdata [30] ), .Z(\AXI4Interconnect/_0328_ ) );
BUF_X1 \AXI4Interconnect/_1628_ ( .A(\io_master_rdata [30] ), .Z(\AXI4Interconnect/_0476_ ) );
BUF_X1 \AXI4Interconnect/_1629_ ( .A(\AXI4Interconnect/_0067_ ), .Z(\_AXI4Interconnect_io_fanIn_0_rdata [30] ) );
BUF_X1 \AXI4Interconnect/_1630_ ( .A(\_CLINT_io_rdata [31] ), .Z(\AXI4Interconnect/_0329_ ) );
BUF_X1 \AXI4Interconnect/_1631_ ( .A(\io_master_rdata [31] ), .Z(\AXI4Interconnect/_0477_ ) );
BUF_X1 \AXI4Interconnect/_1632_ ( .A(\AXI4Interconnect/_0068_ ), .Z(\_AXI4Interconnect_io_fanIn_0_rdata [31] ) );
BUF_X1 \AXI4Interconnect/_1633_ ( .A(\_CLINT_io_bresp [0] ), .Z(\AXI4Interconnect/_0302_ ) );
BUF_X1 \AXI4Interconnect/_1634_ ( .A(\io_master_bresp [0] ), .Z(\AXI4Interconnect/_0450_ ) );
BUF_X1 \AXI4Interconnect/_1635_ ( .A(\AXI4Interconnect/selectedReg ), .Z(\AXI4Interconnect/_0871_ ) );
BUF_X1 \AXI4Interconnect/_1636_ ( .A(\AXI4Interconnect/_0155_ ), .Z(\_AXI4Interconnect_io_fanIn_1_bresp [0] ) );
BUF_X1 \AXI4Interconnect/_1637_ ( .A(\_CLINT_io_bresp [1] ), .Z(\AXI4Interconnect/_0303_ ) );
BUF_X1 \AXI4Interconnect/_1638_ ( .A(\io_master_bresp [1] ), .Z(\AXI4Interconnect/_0451_ ) );
BUF_X1 \AXI4Interconnect/_1639_ ( .A(\AXI4Interconnect/_0156_ ), .Z(\_AXI4Interconnect_io_fanIn_1_bresp [1] ) );
BUF_X1 \AXI4Interconnect/_1640_ ( .A(\AXI4Interconnect/_0191_ ), .Z(\_AXI4Interconnect_io_fanIn_1_rresp [0] ) );
BUF_X1 \AXI4Interconnect/_1641_ ( .A(\AXI4Interconnect/_0192_ ), .Z(\_AXI4Interconnect_io_fanIn_1_rresp [1] ) );
BUF_X1 \AXI4Interconnect/_1642_ ( .A(\AXI4Interconnect/_0158_ ), .Z(\_AXI4Interconnect_io_fanIn_1_rdata [0] ) );
BUF_X1 \AXI4Interconnect/_1643_ ( .A(\AXI4Interconnect/_0169_ ), .Z(\_AXI4Interconnect_io_fanIn_1_rdata [1] ) );
BUF_X1 \AXI4Interconnect/_1644_ ( .A(\AXI4Interconnect/_0180_ ), .Z(\_AXI4Interconnect_io_fanIn_1_rdata [2] ) );
BUF_X1 \AXI4Interconnect/_1645_ ( .A(\AXI4Interconnect/_0183_ ), .Z(\_AXI4Interconnect_io_fanIn_1_rdata [3] ) );
BUF_X1 \AXI4Interconnect/_1646_ ( .A(\AXI4Interconnect/_0184_ ), .Z(\_AXI4Interconnect_io_fanIn_1_rdata [4] ) );
BUF_X1 \AXI4Interconnect/_1647_ ( .A(\AXI4Interconnect/_0185_ ), .Z(\_AXI4Interconnect_io_fanIn_1_rdata [5] ) );
BUF_X1 \AXI4Interconnect/_1648_ ( .A(\AXI4Interconnect/_0186_ ), .Z(\_AXI4Interconnect_io_fanIn_1_rdata [6] ) );
BUF_X1 \AXI4Interconnect/_1649_ ( .A(\AXI4Interconnect/_0187_ ), .Z(\_AXI4Interconnect_io_fanIn_1_rdata [7] ) );
BUF_X1 \AXI4Interconnect/_1650_ ( .A(\AXI4Interconnect/_0188_ ), .Z(\_AXI4Interconnect_io_fanIn_1_rdata [8] ) );
BUF_X1 \AXI4Interconnect/_1651_ ( .A(\AXI4Interconnect/_0189_ ), .Z(\_AXI4Interconnect_io_fanIn_1_rdata [9] ) );
BUF_X1 \AXI4Interconnect/_1652_ ( .A(\AXI4Interconnect/_0159_ ), .Z(\_AXI4Interconnect_io_fanIn_1_rdata [10] ) );
BUF_X1 \AXI4Interconnect/_1653_ ( .A(\AXI4Interconnect/_0160_ ), .Z(\_AXI4Interconnect_io_fanIn_1_rdata [11] ) );
BUF_X1 \AXI4Interconnect/_1654_ ( .A(\AXI4Interconnect/_0161_ ), .Z(\_AXI4Interconnect_io_fanIn_1_rdata [12] ) );
BUF_X1 \AXI4Interconnect/_1655_ ( .A(\AXI4Interconnect/_0162_ ), .Z(\_AXI4Interconnect_io_fanIn_1_rdata [13] ) );
BUF_X1 \AXI4Interconnect/_1656_ ( .A(\AXI4Interconnect/_0163_ ), .Z(\_AXI4Interconnect_io_fanIn_1_rdata [14] ) );
BUF_X1 \AXI4Interconnect/_1657_ ( .A(\AXI4Interconnect/_0164_ ), .Z(\_AXI4Interconnect_io_fanIn_1_rdata [15] ) );
BUF_X1 \AXI4Interconnect/_1658_ ( .A(\AXI4Interconnect/_0165_ ), .Z(\_AXI4Interconnect_io_fanIn_1_rdata [16] ) );
BUF_X1 \AXI4Interconnect/_1659_ ( .A(\AXI4Interconnect/_0166_ ), .Z(\_AXI4Interconnect_io_fanIn_1_rdata [17] ) );
BUF_X1 \AXI4Interconnect/_1660_ ( .A(\AXI4Interconnect/_0167_ ), .Z(\_AXI4Interconnect_io_fanIn_1_rdata [18] ) );
BUF_X1 \AXI4Interconnect/_1661_ ( .A(\AXI4Interconnect/_0168_ ), .Z(\_AXI4Interconnect_io_fanIn_1_rdata [19] ) );
BUF_X1 \AXI4Interconnect/_1662_ ( .A(\AXI4Interconnect/_0170_ ), .Z(\_AXI4Interconnect_io_fanIn_1_rdata [20] ) );
BUF_X1 \AXI4Interconnect/_1663_ ( .A(\AXI4Interconnect/_0171_ ), .Z(\_AXI4Interconnect_io_fanIn_1_rdata [21] ) );
BUF_X1 \AXI4Interconnect/_1664_ ( .A(\AXI4Interconnect/_0172_ ), .Z(\_AXI4Interconnect_io_fanIn_1_rdata [22] ) );
BUF_X1 \AXI4Interconnect/_1665_ ( .A(\AXI4Interconnect/_0173_ ), .Z(\_AXI4Interconnect_io_fanIn_1_rdata [23] ) );
BUF_X1 \AXI4Interconnect/_1666_ ( .A(\AXI4Interconnect/_0174_ ), .Z(\_AXI4Interconnect_io_fanIn_1_rdata [24] ) );
BUF_X1 \AXI4Interconnect/_1667_ ( .A(\AXI4Interconnect/_0175_ ), .Z(\_AXI4Interconnect_io_fanIn_1_rdata [25] ) );
BUF_X1 \AXI4Interconnect/_1668_ ( .A(\AXI4Interconnect/_0176_ ), .Z(\_AXI4Interconnect_io_fanIn_1_rdata [26] ) );
BUF_X1 \AXI4Interconnect/_1669_ ( .A(\AXI4Interconnect/_0177_ ), .Z(\_AXI4Interconnect_io_fanIn_1_rdata [27] ) );
BUF_X1 \AXI4Interconnect/_1670_ ( .A(\AXI4Interconnect/_0178_ ), .Z(\_AXI4Interconnect_io_fanIn_1_rdata [28] ) );
BUF_X1 \AXI4Interconnect/_1671_ ( .A(\AXI4Interconnect/_0179_ ), .Z(\_AXI4Interconnect_io_fanIn_1_rdata [29] ) );
BUF_X1 \AXI4Interconnect/_1672_ ( .A(\AXI4Interconnect/_0181_ ), .Z(\_AXI4Interconnect_io_fanIn_1_rdata [30] ) );
BUF_X1 \AXI4Interconnect/_1673_ ( .A(\AXI4Interconnect/_0182_ ), .Z(\_AXI4Interconnect_io_fanIn_1_rdata [31] ) );
BUF_X1 \AXI4Interconnect/_1674_ ( .A(\AXI4Interconnect/_0001_ ), .Z(\AXI4Interconnect/_0005_ ) );
BUF_X1 \AXI4Interconnect/_1675_ ( .A(\_LSU_io_master_awaddr [0] ), .Z(\AXI4Interconnect/_0117_ ) );
BUF_X1 \AXI4Interconnect/_1676_ ( .A(\AXI4Interconnect/_0267_ ), .Z(\_AXI4Interconnect_io_fanOut_0_awaddr [0] ) );
BUF_X1 \AXI4Interconnect/_1677_ ( .A(\_LSU_io_master_awaddr [1] ), .Z(\AXI4Interconnect/_0128_ ) );
BUF_X1 \AXI4Interconnect/_1678_ ( .A(\AXI4Interconnect/_0278_ ), .Z(\_AXI4Interconnect_io_fanOut_0_awaddr [1] ) );
BUF_X1 \AXI4Interconnect/_1679_ ( .A(\_LSU_io_master_awaddr [2] ), .Z(\AXI4Interconnect/_0139_ ) );
BUF_X1 \AXI4Interconnect/_1680_ ( .A(\AXI4Interconnect/_0289_ ), .Z(\_AXI4Interconnect_io_fanOut_0_awaddr [2] ) );
BUF_X1 \AXI4Interconnect/_1681_ ( .A(\_LSU_io_master_awaddr [3] ), .Z(\AXI4Interconnect/_0142_ ) );
BUF_X1 \AXI4Interconnect/_1682_ ( .A(\AXI4Interconnect/_0292_ ), .Z(\_AXI4Interconnect_io_fanOut_0_awaddr [3] ) );
BUF_X1 \AXI4Interconnect/_1683_ ( .A(\_LSU_io_master_awaddr [4] ), .Z(\AXI4Interconnect/_0143_ ) );
BUF_X1 \AXI4Interconnect/_1684_ ( .A(\AXI4Interconnect/_0293_ ), .Z(\_AXI4Interconnect_io_fanOut_0_awaddr [4] ) );
BUF_X1 \AXI4Interconnect/_1685_ ( .A(\_LSU_io_master_awaddr [5] ), .Z(\AXI4Interconnect/_0144_ ) );
BUF_X1 \AXI4Interconnect/_1686_ ( .A(\AXI4Interconnect/_0294_ ), .Z(\_AXI4Interconnect_io_fanOut_0_awaddr [5] ) );
BUF_X1 \AXI4Interconnect/_1687_ ( .A(\_LSU_io_master_awaddr [6] ), .Z(\AXI4Interconnect/_0145_ ) );
BUF_X1 \AXI4Interconnect/_1688_ ( .A(\AXI4Interconnect/_0295_ ), .Z(\_AXI4Interconnect_io_fanOut_0_awaddr [6] ) );
BUF_X1 \AXI4Interconnect/_1689_ ( .A(\_LSU_io_master_awaddr [7] ), .Z(\AXI4Interconnect/_0146_ ) );
BUF_X1 \AXI4Interconnect/_1690_ ( .A(\AXI4Interconnect/_0296_ ), .Z(\_AXI4Interconnect_io_fanOut_0_awaddr [7] ) );
BUF_X1 \AXI4Interconnect/_1691_ ( .A(\_LSU_io_master_awaddr [8] ), .Z(\AXI4Interconnect/_0147_ ) );
BUF_X1 \AXI4Interconnect/_1692_ ( .A(\AXI4Interconnect/_0297_ ), .Z(\_AXI4Interconnect_io_fanOut_0_awaddr [8] ) );
BUF_X1 \AXI4Interconnect/_1693_ ( .A(\_LSU_io_master_awaddr [9] ), .Z(\AXI4Interconnect/_0148_ ) );
BUF_X1 \AXI4Interconnect/_1694_ ( .A(\AXI4Interconnect/_0298_ ), .Z(\_AXI4Interconnect_io_fanOut_0_awaddr [9] ) );
BUF_X1 \AXI4Interconnect/_1695_ ( .A(\_LSU_io_master_awaddr [10] ), .Z(\AXI4Interconnect/_0118_ ) );
BUF_X1 \AXI4Interconnect/_1696_ ( .A(\AXI4Interconnect/_0268_ ), .Z(\_AXI4Interconnect_io_fanOut_0_awaddr [10] ) );
BUF_X1 \AXI4Interconnect/_1697_ ( .A(\_LSU_io_master_awaddr [11] ), .Z(\AXI4Interconnect/_0119_ ) );
BUF_X1 \AXI4Interconnect/_1698_ ( .A(\AXI4Interconnect/_0269_ ), .Z(\_AXI4Interconnect_io_fanOut_0_awaddr [11] ) );
BUF_X1 \AXI4Interconnect/_1699_ ( .A(\_LSU_io_master_awaddr [12] ), .Z(\AXI4Interconnect/_0120_ ) );
BUF_X1 \AXI4Interconnect/_1700_ ( .A(\AXI4Interconnect/_0270_ ), .Z(\_AXI4Interconnect_io_fanOut_0_awaddr [12] ) );
BUF_X1 \AXI4Interconnect/_1701_ ( .A(\_LSU_io_master_awaddr [13] ), .Z(\AXI4Interconnect/_0121_ ) );
BUF_X1 \AXI4Interconnect/_1702_ ( .A(\AXI4Interconnect/_0271_ ), .Z(\_AXI4Interconnect_io_fanOut_0_awaddr [13] ) );
BUF_X1 \AXI4Interconnect/_1703_ ( .A(\_LSU_io_master_awaddr [14] ), .Z(\AXI4Interconnect/_0122_ ) );
BUF_X1 \AXI4Interconnect/_1704_ ( .A(\AXI4Interconnect/_0272_ ), .Z(\_AXI4Interconnect_io_fanOut_0_awaddr [14] ) );
BUF_X1 \AXI4Interconnect/_1705_ ( .A(\_LSU_io_master_awaddr [15] ), .Z(\AXI4Interconnect/_0123_ ) );
BUF_X1 \AXI4Interconnect/_1706_ ( .A(\AXI4Interconnect/_0273_ ), .Z(\_AXI4Interconnect_io_fanOut_0_awaddr [15] ) );
BUF_X1 \AXI4Interconnect/_1707_ ( .A(\_LSU_io_master_awaddr [16] ), .Z(\AXI4Interconnect/_0124_ ) );
BUF_X1 \AXI4Interconnect/_1708_ ( .A(\AXI4Interconnect/_0274_ ), .Z(\_AXI4Interconnect_io_fanOut_0_awaddr [16] ) );
BUF_X1 \AXI4Interconnect/_1709_ ( .A(\_LSU_io_master_awaddr [17] ), .Z(\AXI4Interconnect/_0125_ ) );
BUF_X1 \AXI4Interconnect/_1710_ ( .A(\AXI4Interconnect/_0275_ ), .Z(\_AXI4Interconnect_io_fanOut_0_awaddr [17] ) );
BUF_X1 \AXI4Interconnect/_1711_ ( .A(\_LSU_io_master_awaddr [18] ), .Z(\AXI4Interconnect/_0126_ ) );
BUF_X1 \AXI4Interconnect/_1712_ ( .A(\AXI4Interconnect/_0276_ ), .Z(\_AXI4Interconnect_io_fanOut_0_awaddr [18] ) );
BUF_X1 \AXI4Interconnect/_1713_ ( .A(\_LSU_io_master_awaddr [19] ), .Z(\AXI4Interconnect/_0127_ ) );
BUF_X1 \AXI4Interconnect/_1714_ ( .A(\AXI4Interconnect/_0277_ ), .Z(\_AXI4Interconnect_io_fanOut_0_awaddr [19] ) );
BUF_X1 \AXI4Interconnect/_1715_ ( .A(\_LSU_io_master_awaddr [20] ), .Z(\AXI4Interconnect/_0129_ ) );
BUF_X1 \AXI4Interconnect/_1716_ ( .A(\AXI4Interconnect/_0279_ ), .Z(\_AXI4Interconnect_io_fanOut_0_awaddr [20] ) );
BUF_X1 \AXI4Interconnect/_1717_ ( .A(\_LSU_io_master_awaddr [21] ), .Z(\AXI4Interconnect/_0130_ ) );
BUF_X1 \AXI4Interconnect/_1718_ ( .A(\AXI4Interconnect/_0280_ ), .Z(\_AXI4Interconnect_io_fanOut_0_awaddr [21] ) );
BUF_X1 \AXI4Interconnect/_1719_ ( .A(\_LSU_io_master_awaddr [22] ), .Z(\AXI4Interconnect/_0131_ ) );
BUF_X1 \AXI4Interconnect/_1720_ ( .A(\AXI4Interconnect/_0281_ ), .Z(\_AXI4Interconnect_io_fanOut_0_awaddr [22] ) );
BUF_X1 \AXI4Interconnect/_1721_ ( .A(\_LSU_io_master_awaddr [23] ), .Z(\AXI4Interconnect/_0132_ ) );
BUF_X1 \AXI4Interconnect/_1722_ ( .A(\AXI4Interconnect/_0282_ ), .Z(\_AXI4Interconnect_io_fanOut_0_awaddr [23] ) );
BUF_X1 \AXI4Interconnect/_1723_ ( .A(\_LSU_io_master_awaddr [24] ), .Z(\AXI4Interconnect/_0133_ ) );
BUF_X1 \AXI4Interconnect/_1724_ ( .A(\AXI4Interconnect/_0283_ ), .Z(\_AXI4Interconnect_io_fanOut_0_awaddr [24] ) );
BUF_X1 \AXI4Interconnect/_1725_ ( .A(\_LSU_io_master_awaddr [25] ), .Z(\AXI4Interconnect/_0134_ ) );
BUF_X1 \AXI4Interconnect/_1726_ ( .A(\AXI4Interconnect/_0284_ ), .Z(\_AXI4Interconnect_io_fanOut_0_awaddr [25] ) );
BUF_X1 \AXI4Interconnect/_1727_ ( .A(\_LSU_io_master_awaddr [26] ), .Z(\AXI4Interconnect/_0135_ ) );
BUF_X1 \AXI4Interconnect/_1728_ ( .A(\AXI4Interconnect/_0285_ ), .Z(\_AXI4Interconnect_io_fanOut_0_awaddr [26] ) );
BUF_X1 \AXI4Interconnect/_1729_ ( .A(\_LSU_io_master_awaddr [27] ), .Z(\AXI4Interconnect/_0136_ ) );
BUF_X1 \AXI4Interconnect/_1730_ ( .A(\AXI4Interconnect/_0286_ ), .Z(\_AXI4Interconnect_io_fanOut_0_awaddr [27] ) );
BUF_X1 \AXI4Interconnect/_1731_ ( .A(\_LSU_io_master_awaddr [28] ), .Z(\AXI4Interconnect/_0137_ ) );
BUF_X1 \AXI4Interconnect/_1732_ ( .A(\AXI4Interconnect/_0287_ ), .Z(\_AXI4Interconnect_io_fanOut_0_awaddr [28] ) );
BUF_X1 \AXI4Interconnect/_1733_ ( .A(\_LSU_io_master_awaddr [29] ), .Z(\AXI4Interconnect/_0138_ ) );
BUF_X1 \AXI4Interconnect/_1734_ ( .A(\AXI4Interconnect/_0288_ ), .Z(\_AXI4Interconnect_io_fanOut_0_awaddr [29] ) );
BUF_X1 \AXI4Interconnect/_1735_ ( .A(\_LSU_io_master_awaddr [30] ), .Z(\AXI4Interconnect/_0140_ ) );
BUF_X1 \AXI4Interconnect/_1736_ ( .A(\AXI4Interconnect/_0290_ ), .Z(\_AXI4Interconnect_io_fanOut_0_awaddr [30] ) );
BUF_X1 \AXI4Interconnect/_1737_ ( .A(\_LSU_io_master_awaddr [31] ), .Z(\AXI4Interconnect/_0141_ ) );
BUF_X1 \AXI4Interconnect/_1738_ ( .A(\AXI4Interconnect/_0291_ ), .Z(\_AXI4Interconnect_io_fanOut_0_awaddr [31] ) );
BUF_X1 \AXI4Interconnect/_1739_ ( .A(\_LSU_io_master_wdata [0] ), .Z(\AXI4Interconnect/_0194_ ) );
BUF_X1 \AXI4Interconnect/_1740_ ( .A(\AXI4Interconnect/_0341_ ), .Z(\_AXI4Interconnect_io_fanOut_0_wdata [0] ) );
BUF_X1 \AXI4Interconnect/_1741_ ( .A(\_LSU_io_master_wdata [1] ), .Z(\AXI4Interconnect/_0205_ ) );
BUF_X1 \AXI4Interconnect/_1742_ ( .A(\AXI4Interconnect/_0352_ ), .Z(\_AXI4Interconnect_io_fanOut_0_wdata [1] ) );
BUF_X1 \AXI4Interconnect/_1743_ ( .A(\_LSU_io_master_wdata [2] ), .Z(\AXI4Interconnect/_0216_ ) );
BUF_X1 \AXI4Interconnect/_1744_ ( .A(\AXI4Interconnect/_0363_ ), .Z(\_AXI4Interconnect_io_fanOut_0_wdata [2] ) );
BUF_X1 \AXI4Interconnect/_1745_ ( .A(\_LSU_io_master_wdata [3] ), .Z(\AXI4Interconnect/_0219_ ) );
BUF_X1 \AXI4Interconnect/_1746_ ( .A(\AXI4Interconnect/_0366_ ), .Z(\_AXI4Interconnect_io_fanOut_0_wdata [3] ) );
BUF_X1 \AXI4Interconnect/_1747_ ( .A(\_LSU_io_master_wdata [4] ), .Z(\AXI4Interconnect/_0220_ ) );
BUF_X1 \AXI4Interconnect/_1748_ ( .A(\AXI4Interconnect/_0367_ ), .Z(\_AXI4Interconnect_io_fanOut_0_wdata [4] ) );
BUF_X1 \AXI4Interconnect/_1749_ ( .A(\_LSU_io_master_wdata [5] ), .Z(\AXI4Interconnect/_0221_ ) );
BUF_X1 \AXI4Interconnect/_1750_ ( .A(\AXI4Interconnect/_0368_ ), .Z(\_AXI4Interconnect_io_fanOut_0_wdata [5] ) );
BUF_X1 \AXI4Interconnect/_1751_ ( .A(\_LSU_io_master_wdata [6] ), .Z(\AXI4Interconnect/_0222_ ) );
BUF_X1 \AXI4Interconnect/_1752_ ( .A(\AXI4Interconnect/_0369_ ), .Z(\_AXI4Interconnect_io_fanOut_0_wdata [6] ) );
BUF_X1 \AXI4Interconnect/_1753_ ( .A(\_LSU_io_master_wdata [7] ), .Z(\AXI4Interconnect/_0223_ ) );
BUF_X1 \AXI4Interconnect/_1754_ ( .A(\AXI4Interconnect/_0370_ ), .Z(\_AXI4Interconnect_io_fanOut_0_wdata [7] ) );
BUF_X1 \AXI4Interconnect/_1755_ ( .A(\_LSU_io_master_wdata [8] ), .Z(\AXI4Interconnect/_0224_ ) );
BUF_X1 \AXI4Interconnect/_1756_ ( .A(\AXI4Interconnect/_0371_ ), .Z(\_AXI4Interconnect_io_fanOut_0_wdata [8] ) );
BUF_X1 \AXI4Interconnect/_1757_ ( .A(\_LSU_io_master_wdata [9] ), .Z(\AXI4Interconnect/_0225_ ) );
BUF_X1 \AXI4Interconnect/_1758_ ( .A(\AXI4Interconnect/_0372_ ), .Z(\_AXI4Interconnect_io_fanOut_0_wdata [9] ) );
BUF_X1 \AXI4Interconnect/_1759_ ( .A(\_LSU_io_master_wdata [10] ), .Z(\AXI4Interconnect/_0195_ ) );
BUF_X1 \AXI4Interconnect/_1760_ ( .A(\AXI4Interconnect/_0342_ ), .Z(\_AXI4Interconnect_io_fanOut_0_wdata [10] ) );
BUF_X1 \AXI4Interconnect/_1761_ ( .A(\_LSU_io_master_wdata [11] ), .Z(\AXI4Interconnect/_0196_ ) );
BUF_X1 \AXI4Interconnect/_1762_ ( .A(\AXI4Interconnect/_0343_ ), .Z(\_AXI4Interconnect_io_fanOut_0_wdata [11] ) );
BUF_X1 \AXI4Interconnect/_1763_ ( .A(\_LSU_io_master_wdata [12] ), .Z(\AXI4Interconnect/_0197_ ) );
BUF_X1 \AXI4Interconnect/_1764_ ( .A(\AXI4Interconnect/_0344_ ), .Z(\_AXI4Interconnect_io_fanOut_0_wdata [12] ) );
BUF_X1 \AXI4Interconnect/_1765_ ( .A(\_LSU_io_master_wdata [13] ), .Z(\AXI4Interconnect/_0198_ ) );
BUF_X1 \AXI4Interconnect/_1766_ ( .A(\AXI4Interconnect/_0345_ ), .Z(\_AXI4Interconnect_io_fanOut_0_wdata [13] ) );
BUF_X1 \AXI4Interconnect/_1767_ ( .A(\_LSU_io_master_wdata [14] ), .Z(\AXI4Interconnect/_0199_ ) );
BUF_X1 \AXI4Interconnect/_1768_ ( .A(\AXI4Interconnect/_0346_ ), .Z(\_AXI4Interconnect_io_fanOut_0_wdata [14] ) );
BUF_X1 \AXI4Interconnect/_1769_ ( .A(\_LSU_io_master_wdata [15] ), .Z(\AXI4Interconnect/_0200_ ) );
BUF_X1 \AXI4Interconnect/_1770_ ( .A(\AXI4Interconnect/_0347_ ), .Z(\_AXI4Interconnect_io_fanOut_0_wdata [15] ) );
BUF_X1 \AXI4Interconnect/_1771_ ( .A(\_LSU_io_master_wdata [16] ), .Z(\AXI4Interconnect/_0201_ ) );
BUF_X1 \AXI4Interconnect/_1772_ ( .A(\AXI4Interconnect/_0348_ ), .Z(\_AXI4Interconnect_io_fanOut_0_wdata [16] ) );
BUF_X1 \AXI4Interconnect/_1773_ ( .A(\_LSU_io_master_wdata [17] ), .Z(\AXI4Interconnect/_0202_ ) );
BUF_X1 \AXI4Interconnect/_1774_ ( .A(\AXI4Interconnect/_0349_ ), .Z(\_AXI4Interconnect_io_fanOut_0_wdata [17] ) );
BUF_X1 \AXI4Interconnect/_1775_ ( .A(\_LSU_io_master_wdata [18] ), .Z(\AXI4Interconnect/_0203_ ) );
BUF_X1 \AXI4Interconnect/_1776_ ( .A(\AXI4Interconnect/_0350_ ), .Z(\_AXI4Interconnect_io_fanOut_0_wdata [18] ) );
BUF_X1 \AXI4Interconnect/_1777_ ( .A(\_LSU_io_master_wdata [19] ), .Z(\AXI4Interconnect/_0204_ ) );
BUF_X1 \AXI4Interconnect/_1778_ ( .A(\AXI4Interconnect/_0351_ ), .Z(\_AXI4Interconnect_io_fanOut_0_wdata [19] ) );
BUF_X1 \AXI4Interconnect/_1779_ ( .A(\_LSU_io_master_wdata [20] ), .Z(\AXI4Interconnect/_0206_ ) );
BUF_X1 \AXI4Interconnect/_1780_ ( .A(\AXI4Interconnect/_0353_ ), .Z(\_AXI4Interconnect_io_fanOut_0_wdata [20] ) );
BUF_X1 \AXI4Interconnect/_1781_ ( .A(\_LSU_io_master_wdata [21] ), .Z(\AXI4Interconnect/_0207_ ) );
BUF_X1 \AXI4Interconnect/_1782_ ( .A(\AXI4Interconnect/_0354_ ), .Z(\_AXI4Interconnect_io_fanOut_0_wdata [21] ) );
BUF_X1 \AXI4Interconnect/_1783_ ( .A(\_LSU_io_master_wdata [22] ), .Z(\AXI4Interconnect/_0208_ ) );
BUF_X1 \AXI4Interconnect/_1784_ ( .A(\AXI4Interconnect/_0355_ ), .Z(\_AXI4Interconnect_io_fanOut_0_wdata [22] ) );
BUF_X1 \AXI4Interconnect/_1785_ ( .A(\_LSU_io_master_wdata [23] ), .Z(\AXI4Interconnect/_0209_ ) );
BUF_X1 \AXI4Interconnect/_1786_ ( .A(\AXI4Interconnect/_0356_ ), .Z(\_AXI4Interconnect_io_fanOut_0_wdata [23] ) );
BUF_X1 \AXI4Interconnect/_1787_ ( .A(\_LSU_io_master_wdata [24] ), .Z(\AXI4Interconnect/_0210_ ) );
BUF_X1 \AXI4Interconnect/_1788_ ( .A(\AXI4Interconnect/_0357_ ), .Z(\_AXI4Interconnect_io_fanOut_0_wdata [24] ) );
BUF_X1 \AXI4Interconnect/_1789_ ( .A(\_LSU_io_master_wdata [25] ), .Z(\AXI4Interconnect/_0211_ ) );
BUF_X1 \AXI4Interconnect/_1790_ ( .A(\AXI4Interconnect/_0358_ ), .Z(\_AXI4Interconnect_io_fanOut_0_wdata [25] ) );
BUF_X1 \AXI4Interconnect/_1791_ ( .A(\_LSU_io_master_wdata [26] ), .Z(\AXI4Interconnect/_0212_ ) );
BUF_X1 \AXI4Interconnect/_1792_ ( .A(\AXI4Interconnect/_0359_ ), .Z(\_AXI4Interconnect_io_fanOut_0_wdata [26] ) );
BUF_X1 \AXI4Interconnect/_1793_ ( .A(\_LSU_io_master_wdata [27] ), .Z(\AXI4Interconnect/_0213_ ) );
BUF_X1 \AXI4Interconnect/_1794_ ( .A(\AXI4Interconnect/_0360_ ), .Z(\_AXI4Interconnect_io_fanOut_0_wdata [27] ) );
BUF_X1 \AXI4Interconnect/_1795_ ( .A(\_LSU_io_master_wdata [28] ), .Z(\AXI4Interconnect/_0214_ ) );
BUF_X1 \AXI4Interconnect/_1796_ ( .A(\AXI4Interconnect/_0361_ ), .Z(\_AXI4Interconnect_io_fanOut_0_wdata [28] ) );
BUF_X1 \AXI4Interconnect/_1797_ ( .A(\_LSU_io_master_wdata [29] ), .Z(\AXI4Interconnect/_0215_ ) );
BUF_X1 \AXI4Interconnect/_1798_ ( .A(\AXI4Interconnect/_0362_ ), .Z(\_AXI4Interconnect_io_fanOut_0_wdata [29] ) );
BUF_X1 \AXI4Interconnect/_1799_ ( .A(\_LSU_io_master_wdata [30] ), .Z(\AXI4Interconnect/_0217_ ) );
BUF_X1 \AXI4Interconnect/_1800_ ( .A(\AXI4Interconnect/_0364_ ), .Z(\_AXI4Interconnect_io_fanOut_0_wdata [30] ) );
BUF_X1 \AXI4Interconnect/_1801_ ( .A(\_LSU_io_master_wdata [31] ), .Z(\AXI4Interconnect/_0218_ ) );
BUF_X1 \AXI4Interconnect/_1802_ ( .A(\AXI4Interconnect/_0365_ ), .Z(\_AXI4Interconnect_io_fanOut_0_wdata [31] ) );
BUF_X1 \AXI4Interconnect/_1803_ ( .A(\_IFU_io_master_araddr [0] ), .Z(\AXI4Interconnect/_0010_ ) );
BUF_X1 \AXI4Interconnect/_1804_ ( .A(\_LSU_io_master_araddr [0] ), .Z(\AXI4Interconnect/_0080_ ) );
BUF_X1 \AXI4Interconnect/_1805_ ( .A(\AXI4Interconnect/_0233_ ), .Z(\_AXI4Interconnect_io_fanOut_0_araddr [0] ) );
BUF_X1 \AXI4Interconnect/_1806_ ( .A(\_IFU_io_master_araddr [1] ), .Z(\AXI4Interconnect/_0021_ ) );
BUF_X1 \AXI4Interconnect/_1807_ ( .A(\_LSU_io_master_araddr [1] ), .Z(\AXI4Interconnect/_0091_ ) );
BUF_X1 \AXI4Interconnect/_1808_ ( .A(\AXI4Interconnect/_0244_ ), .Z(\_AXI4Interconnect_io_fanOut_0_araddr [1] ) );
BUF_X1 \AXI4Interconnect/_1809_ ( .A(\_IFU_io_master_araddr [2] ), .Z(\AXI4Interconnect/_0032_ ) );
BUF_X1 \AXI4Interconnect/_1810_ ( .A(\_LSU_io_master_araddr [2] ), .Z(\AXI4Interconnect/_0102_ ) );
BUF_X1 \AXI4Interconnect/_1811_ ( .A(\AXI4Interconnect/_0255_ ), .Z(\_AXI4Interconnect_io_fanOut_0_araddr [2] ) );
BUF_X1 \AXI4Interconnect/_1812_ ( .A(\_IFU_io_master_araddr [3] ), .Z(\AXI4Interconnect/_0035_ ) );
BUF_X1 \AXI4Interconnect/_1813_ ( .A(\_LSU_io_master_araddr [3] ), .Z(\AXI4Interconnect/_0105_ ) );
BUF_X1 \AXI4Interconnect/_1814_ ( .A(\AXI4Interconnect/_0258_ ), .Z(\_AXI4Interconnect_io_fanOut_0_araddr [3] ) );
BUF_X1 \AXI4Interconnect/_1815_ ( .A(\_IFU_io_master_araddr [4] ), .Z(\AXI4Interconnect/_0036_ ) );
BUF_X1 \AXI4Interconnect/_1816_ ( .A(\_LSU_io_master_araddr [4] ), .Z(\AXI4Interconnect/_0106_ ) );
BUF_X1 \AXI4Interconnect/_1817_ ( .A(\AXI4Interconnect/_0259_ ), .Z(\_AXI4Interconnect_io_fanOut_0_araddr [4] ) );
BUF_X1 \AXI4Interconnect/_1818_ ( .A(\_IFU_io_master_araddr [5] ), .Z(\AXI4Interconnect/_0037_ ) );
BUF_X1 \AXI4Interconnect/_1819_ ( .A(\_LSU_io_master_araddr [5] ), .Z(\AXI4Interconnect/_0107_ ) );
BUF_X1 \AXI4Interconnect/_1820_ ( .A(\AXI4Interconnect/_0260_ ), .Z(\_AXI4Interconnect_io_fanOut_0_araddr [5] ) );
BUF_X1 \AXI4Interconnect/_1821_ ( .A(\_IFU_io_master_araddr [6] ), .Z(\AXI4Interconnect/_0038_ ) );
BUF_X1 \AXI4Interconnect/_1822_ ( .A(\_LSU_io_master_araddr [6] ), .Z(\AXI4Interconnect/_0108_ ) );
BUF_X1 \AXI4Interconnect/_1823_ ( .A(\AXI4Interconnect/_0261_ ), .Z(\_AXI4Interconnect_io_fanOut_0_araddr [6] ) );
BUF_X1 \AXI4Interconnect/_1824_ ( .A(\_IFU_io_master_araddr [7] ), .Z(\AXI4Interconnect/_0039_ ) );
BUF_X1 \AXI4Interconnect/_1825_ ( .A(\_LSU_io_master_araddr [7] ), .Z(\AXI4Interconnect/_0109_ ) );
BUF_X1 \AXI4Interconnect/_1826_ ( .A(\AXI4Interconnect/_0262_ ), .Z(\_AXI4Interconnect_io_fanOut_0_araddr [7] ) );
BUF_X1 \AXI4Interconnect/_1827_ ( .A(\_IFU_io_master_araddr [8] ), .Z(\AXI4Interconnect/_0040_ ) );
BUF_X1 \AXI4Interconnect/_1828_ ( .A(\_LSU_io_master_araddr [8] ), .Z(\AXI4Interconnect/_0110_ ) );
BUF_X1 \AXI4Interconnect/_1829_ ( .A(\AXI4Interconnect/_0263_ ), .Z(\_AXI4Interconnect_io_fanOut_0_araddr [8] ) );
BUF_X1 \AXI4Interconnect/_1830_ ( .A(\_IFU_io_master_araddr [9] ), .Z(\AXI4Interconnect/_0041_ ) );
BUF_X1 \AXI4Interconnect/_1831_ ( .A(\_LSU_io_master_araddr [9] ), .Z(\AXI4Interconnect/_0111_ ) );
BUF_X1 \AXI4Interconnect/_1832_ ( .A(\AXI4Interconnect/_0264_ ), .Z(\_AXI4Interconnect_io_fanOut_0_araddr [9] ) );
BUF_X1 \AXI4Interconnect/_1833_ ( .A(\_IFU_io_master_araddr [10] ), .Z(\AXI4Interconnect/_0011_ ) );
BUF_X1 \AXI4Interconnect/_1834_ ( .A(\_LSU_io_master_araddr [10] ), .Z(\AXI4Interconnect/_0081_ ) );
BUF_X1 \AXI4Interconnect/_1835_ ( .A(\AXI4Interconnect/_0234_ ), .Z(\_AXI4Interconnect_io_fanOut_0_araddr [10] ) );
BUF_X1 \AXI4Interconnect/_1836_ ( .A(\_IFU_io_master_araddr [11] ), .Z(\AXI4Interconnect/_0012_ ) );
BUF_X1 \AXI4Interconnect/_1837_ ( .A(\_LSU_io_master_araddr [11] ), .Z(\AXI4Interconnect/_0082_ ) );
BUF_X1 \AXI4Interconnect/_1838_ ( .A(\AXI4Interconnect/_0235_ ), .Z(\_AXI4Interconnect_io_fanOut_0_araddr [11] ) );
BUF_X1 \AXI4Interconnect/_1839_ ( .A(\_IFU_io_master_araddr [12] ), .Z(\AXI4Interconnect/_0013_ ) );
BUF_X1 \AXI4Interconnect/_1840_ ( .A(\_LSU_io_master_araddr [12] ), .Z(\AXI4Interconnect/_0083_ ) );
BUF_X1 \AXI4Interconnect/_1841_ ( .A(\AXI4Interconnect/_0236_ ), .Z(\_AXI4Interconnect_io_fanOut_0_araddr [12] ) );
BUF_X1 \AXI4Interconnect/_1842_ ( .A(\_IFU_io_master_araddr [13] ), .Z(\AXI4Interconnect/_0014_ ) );
BUF_X1 \AXI4Interconnect/_1843_ ( .A(\_LSU_io_master_araddr [13] ), .Z(\AXI4Interconnect/_0084_ ) );
BUF_X1 \AXI4Interconnect/_1844_ ( .A(\AXI4Interconnect/_0237_ ), .Z(\_AXI4Interconnect_io_fanOut_0_araddr [13] ) );
BUF_X1 \AXI4Interconnect/_1845_ ( .A(\_IFU_io_master_araddr [14] ), .Z(\AXI4Interconnect/_0015_ ) );
BUF_X1 \AXI4Interconnect/_1846_ ( .A(\_LSU_io_master_araddr [14] ), .Z(\AXI4Interconnect/_0085_ ) );
BUF_X1 \AXI4Interconnect/_1847_ ( .A(\AXI4Interconnect/_0238_ ), .Z(\_AXI4Interconnect_io_fanOut_0_araddr [14] ) );
BUF_X1 \AXI4Interconnect/_1848_ ( .A(\_IFU_io_master_araddr [15] ), .Z(\AXI4Interconnect/_0016_ ) );
BUF_X1 \AXI4Interconnect/_1849_ ( .A(\_LSU_io_master_araddr [15] ), .Z(\AXI4Interconnect/_0086_ ) );
BUF_X1 \AXI4Interconnect/_1850_ ( .A(\AXI4Interconnect/_0239_ ), .Z(\_AXI4Interconnect_io_fanOut_0_araddr [15] ) );
BUF_X1 \AXI4Interconnect/_1851_ ( .A(\_IFU_io_master_araddr [16] ), .Z(\AXI4Interconnect/_0017_ ) );
BUF_X1 \AXI4Interconnect/_1852_ ( .A(\_LSU_io_master_araddr [16] ), .Z(\AXI4Interconnect/_0087_ ) );
BUF_X1 \AXI4Interconnect/_1853_ ( .A(\AXI4Interconnect/_0240_ ), .Z(\_AXI4Interconnect_io_fanOut_0_araddr [16] ) );
BUF_X1 \AXI4Interconnect/_1854_ ( .A(\_IFU_io_master_araddr [17] ), .Z(\AXI4Interconnect/_0018_ ) );
BUF_X1 \AXI4Interconnect/_1855_ ( .A(\_LSU_io_master_araddr [17] ), .Z(\AXI4Interconnect/_0088_ ) );
BUF_X1 \AXI4Interconnect/_1856_ ( .A(\AXI4Interconnect/_0241_ ), .Z(\_AXI4Interconnect_io_fanOut_0_araddr [17] ) );
BUF_X1 \AXI4Interconnect/_1857_ ( .A(\_IFU_io_master_araddr [18] ), .Z(\AXI4Interconnect/_0019_ ) );
BUF_X1 \AXI4Interconnect/_1858_ ( .A(\_LSU_io_master_araddr [18] ), .Z(\AXI4Interconnect/_0089_ ) );
BUF_X1 \AXI4Interconnect/_1859_ ( .A(\AXI4Interconnect/_0242_ ), .Z(\_AXI4Interconnect_io_fanOut_0_araddr [18] ) );
BUF_X1 \AXI4Interconnect/_1860_ ( .A(\_IFU_io_master_araddr [19] ), .Z(\AXI4Interconnect/_0020_ ) );
BUF_X1 \AXI4Interconnect/_1861_ ( .A(\_LSU_io_master_araddr [19] ), .Z(\AXI4Interconnect/_0090_ ) );
BUF_X1 \AXI4Interconnect/_1862_ ( .A(\AXI4Interconnect/_0243_ ), .Z(\_AXI4Interconnect_io_fanOut_0_araddr [19] ) );
BUF_X1 \AXI4Interconnect/_1863_ ( .A(\_IFU_io_master_araddr [20] ), .Z(\AXI4Interconnect/_0022_ ) );
BUF_X1 \AXI4Interconnect/_1864_ ( .A(\_LSU_io_master_araddr [20] ), .Z(\AXI4Interconnect/_0092_ ) );
BUF_X1 \AXI4Interconnect/_1865_ ( .A(\AXI4Interconnect/_0245_ ), .Z(\_AXI4Interconnect_io_fanOut_0_araddr [20] ) );
BUF_X1 \AXI4Interconnect/_1866_ ( .A(\_IFU_io_master_araddr [21] ), .Z(\AXI4Interconnect/_0023_ ) );
BUF_X1 \AXI4Interconnect/_1867_ ( .A(\_LSU_io_master_araddr [21] ), .Z(\AXI4Interconnect/_0093_ ) );
BUF_X1 \AXI4Interconnect/_1868_ ( .A(\AXI4Interconnect/_0246_ ), .Z(\_AXI4Interconnect_io_fanOut_0_araddr [21] ) );
BUF_X1 \AXI4Interconnect/_1869_ ( .A(\_IFU_io_master_araddr [22] ), .Z(\AXI4Interconnect/_0024_ ) );
BUF_X1 \AXI4Interconnect/_1870_ ( .A(\_LSU_io_master_araddr [22] ), .Z(\AXI4Interconnect/_0094_ ) );
BUF_X1 \AXI4Interconnect/_1871_ ( .A(\AXI4Interconnect/_0247_ ), .Z(\_AXI4Interconnect_io_fanOut_0_araddr [22] ) );
BUF_X1 \AXI4Interconnect/_1872_ ( .A(\_IFU_io_master_araddr [23] ), .Z(\AXI4Interconnect/_0025_ ) );
BUF_X1 \AXI4Interconnect/_1873_ ( .A(\_LSU_io_master_araddr [23] ), .Z(\AXI4Interconnect/_0095_ ) );
BUF_X1 \AXI4Interconnect/_1874_ ( .A(\AXI4Interconnect/_0248_ ), .Z(\_AXI4Interconnect_io_fanOut_0_araddr [23] ) );
BUF_X1 \AXI4Interconnect/_1875_ ( .A(\_IFU_io_master_araddr [24] ), .Z(\AXI4Interconnect/_0026_ ) );
BUF_X1 \AXI4Interconnect/_1876_ ( .A(\_LSU_io_master_araddr [24] ), .Z(\AXI4Interconnect/_0096_ ) );
BUF_X1 \AXI4Interconnect/_1877_ ( .A(\AXI4Interconnect/_0249_ ), .Z(\_AXI4Interconnect_io_fanOut_0_araddr [24] ) );
BUF_X1 \AXI4Interconnect/_1878_ ( .A(\_IFU_io_master_araddr [25] ), .Z(\AXI4Interconnect/_0027_ ) );
BUF_X1 \AXI4Interconnect/_1879_ ( .A(\_LSU_io_master_araddr [25] ), .Z(\AXI4Interconnect/_0097_ ) );
BUF_X1 \AXI4Interconnect/_1880_ ( .A(\AXI4Interconnect/_0250_ ), .Z(\_AXI4Interconnect_io_fanOut_0_araddr [25] ) );
BUF_X1 \AXI4Interconnect/_1881_ ( .A(\_IFU_io_master_araddr [26] ), .Z(\AXI4Interconnect/_0028_ ) );
BUF_X1 \AXI4Interconnect/_1882_ ( .A(\_LSU_io_master_araddr [26] ), .Z(\AXI4Interconnect/_0098_ ) );
BUF_X1 \AXI4Interconnect/_1883_ ( .A(\AXI4Interconnect/_0251_ ), .Z(\_AXI4Interconnect_io_fanOut_0_araddr [26] ) );
BUF_X1 \AXI4Interconnect/_1884_ ( .A(\_IFU_io_master_araddr [27] ), .Z(\AXI4Interconnect/_0029_ ) );
BUF_X1 \AXI4Interconnect/_1885_ ( .A(\_LSU_io_master_araddr [27] ), .Z(\AXI4Interconnect/_0099_ ) );
BUF_X1 \AXI4Interconnect/_1886_ ( .A(\AXI4Interconnect/_0252_ ), .Z(\_AXI4Interconnect_io_fanOut_0_araddr [27] ) );
BUF_X1 \AXI4Interconnect/_1887_ ( .A(\_IFU_io_master_araddr [28] ), .Z(\AXI4Interconnect/_0030_ ) );
BUF_X1 \AXI4Interconnect/_1888_ ( .A(\_LSU_io_master_araddr [28] ), .Z(\AXI4Interconnect/_0100_ ) );
BUF_X1 \AXI4Interconnect/_1889_ ( .A(\AXI4Interconnect/_0253_ ), .Z(\_AXI4Interconnect_io_fanOut_0_araddr [28] ) );
BUF_X1 \AXI4Interconnect/_1890_ ( .A(\_IFU_io_master_araddr [29] ), .Z(\AXI4Interconnect/_0031_ ) );
BUF_X1 \AXI4Interconnect/_1891_ ( .A(\_LSU_io_master_araddr [29] ), .Z(\AXI4Interconnect/_0101_ ) );
BUF_X1 \AXI4Interconnect/_1892_ ( .A(\AXI4Interconnect/_0254_ ), .Z(\_AXI4Interconnect_io_fanOut_0_araddr [29] ) );
BUF_X1 \AXI4Interconnect/_1893_ ( .A(\_IFU_io_master_araddr [30] ), .Z(\AXI4Interconnect/_0033_ ) );
BUF_X1 \AXI4Interconnect/_1894_ ( .A(\_LSU_io_master_araddr [30] ), .Z(\AXI4Interconnect/_0103_ ) );
BUF_X1 \AXI4Interconnect/_1895_ ( .A(\AXI4Interconnect/_0256_ ), .Z(\_AXI4Interconnect_io_fanOut_0_araddr [30] ) );
BUF_X1 \AXI4Interconnect/_1896_ ( .A(\_IFU_io_master_araddr [31] ), .Z(\AXI4Interconnect/_0034_ ) );
BUF_X1 \AXI4Interconnect/_1897_ ( .A(\_LSU_io_master_araddr [31] ), .Z(\AXI4Interconnect/_0104_ ) );
BUF_X1 \AXI4Interconnect/_1898_ ( .A(\AXI4Interconnect/_0257_ ), .Z(\_AXI4Interconnect_io_fanOut_0_araddr [31] ) );
BUF_X1 \AXI4Interconnect/_1899_ ( .A(\AXI4Interconnect/_0002_ ), .Z(\AXI4Interconnect/_GEN_13 ) );
BUF_X1 \AXI4Interconnect/_1900_ ( .A(\AXI4Interconnect/_0003_ ), .Z(\AXI4Interconnect/_GEN_14 ) );
BUF_X1 \AXI4Interconnect/_1901_ ( .A(\AXI4Interconnect/_0412_ ), .Z(\io_master_awaddr [0] ) );
BUF_X1 \AXI4Interconnect/_1902_ ( .A(\AXI4Interconnect/_0423_ ), .Z(\io_master_awaddr [1] ) );
BUF_X1 \AXI4Interconnect/_1903_ ( .A(\AXI4Interconnect/_0434_ ), .Z(\io_master_awaddr [2] ) );
BUF_X1 \AXI4Interconnect/_1904_ ( .A(\AXI4Interconnect/_0437_ ), .Z(\io_master_awaddr [3] ) );
BUF_X1 \AXI4Interconnect/_1905_ ( .A(\AXI4Interconnect/_0438_ ), .Z(\io_master_awaddr [4] ) );
BUF_X1 \AXI4Interconnect/_1906_ ( .A(\AXI4Interconnect/_0439_ ), .Z(\io_master_awaddr [5] ) );
BUF_X1 \AXI4Interconnect/_1907_ ( .A(\AXI4Interconnect/_0440_ ), .Z(\io_master_awaddr [6] ) );
BUF_X1 \AXI4Interconnect/_1908_ ( .A(\AXI4Interconnect/_0441_ ), .Z(\io_master_awaddr [7] ) );
BUF_X1 \AXI4Interconnect/_1909_ ( .A(\AXI4Interconnect/_0442_ ), .Z(\io_master_awaddr [8] ) );
BUF_X1 \AXI4Interconnect/_1910_ ( .A(\AXI4Interconnect/_0443_ ), .Z(\io_master_awaddr [9] ) );
BUF_X1 \AXI4Interconnect/_1911_ ( .A(\AXI4Interconnect/_0413_ ), .Z(\io_master_awaddr [10] ) );
BUF_X1 \AXI4Interconnect/_1912_ ( .A(\AXI4Interconnect/_0414_ ), .Z(\io_master_awaddr [11] ) );
BUF_X1 \AXI4Interconnect/_1913_ ( .A(\AXI4Interconnect/_0415_ ), .Z(\io_master_awaddr [12] ) );
BUF_X1 \AXI4Interconnect/_1914_ ( .A(\AXI4Interconnect/_0416_ ), .Z(\io_master_awaddr [13] ) );
BUF_X1 \AXI4Interconnect/_1915_ ( .A(\AXI4Interconnect/_0417_ ), .Z(\io_master_awaddr [14] ) );
BUF_X1 \AXI4Interconnect/_1916_ ( .A(\AXI4Interconnect/_0418_ ), .Z(\io_master_awaddr [15] ) );
BUF_X1 \AXI4Interconnect/_1917_ ( .A(\AXI4Interconnect/_0419_ ), .Z(\io_master_awaddr [16] ) );
BUF_X1 \AXI4Interconnect/_1918_ ( .A(\AXI4Interconnect/_0420_ ), .Z(\io_master_awaddr [17] ) );
BUF_X1 \AXI4Interconnect/_1919_ ( .A(\AXI4Interconnect/_0421_ ), .Z(\io_master_awaddr [18] ) );
BUF_X1 \AXI4Interconnect/_1920_ ( .A(\AXI4Interconnect/_0422_ ), .Z(\io_master_awaddr [19] ) );
BUF_X1 \AXI4Interconnect/_1921_ ( .A(\AXI4Interconnect/_0424_ ), .Z(\io_master_awaddr [20] ) );
BUF_X1 \AXI4Interconnect/_1922_ ( .A(\AXI4Interconnect/_0425_ ), .Z(\io_master_awaddr [21] ) );
BUF_X1 \AXI4Interconnect/_1923_ ( .A(\AXI4Interconnect/_0426_ ), .Z(\io_master_awaddr [22] ) );
BUF_X1 \AXI4Interconnect/_1924_ ( .A(\AXI4Interconnect/_0427_ ), .Z(\io_master_awaddr [23] ) );
BUF_X1 \AXI4Interconnect/_1925_ ( .A(\AXI4Interconnect/_0428_ ), .Z(\io_master_awaddr [24] ) );
BUF_X1 \AXI4Interconnect/_1926_ ( .A(\AXI4Interconnect/_0429_ ), .Z(\io_master_awaddr [25] ) );
BUF_X1 \AXI4Interconnect/_1927_ ( .A(\AXI4Interconnect/_0430_ ), .Z(\io_master_awaddr [26] ) );
BUF_X1 \AXI4Interconnect/_1928_ ( .A(\AXI4Interconnect/_0431_ ), .Z(\io_master_awaddr [27] ) );
BUF_X1 \AXI4Interconnect/_1929_ ( .A(\AXI4Interconnect/_0432_ ), .Z(\io_master_awaddr [28] ) );
BUF_X1 \AXI4Interconnect/_1930_ ( .A(\AXI4Interconnect/_0433_ ), .Z(\io_master_awaddr [29] ) );
BUF_X1 \AXI4Interconnect/_1931_ ( .A(\AXI4Interconnect/_0435_ ), .Z(\io_master_awaddr [30] ) );
BUF_X1 \AXI4Interconnect/_1932_ ( .A(\AXI4Interconnect/_0436_ ), .Z(\io_master_awaddr [31] ) );
BUF_X1 \AXI4Interconnect/_1933_ ( .A(\AXI4Interconnect/_0489_ ), .Z(\io_master_wdata [0] ) );
BUF_X1 \AXI4Interconnect/_1934_ ( .A(\AXI4Interconnect/_0500_ ), .Z(\io_master_wdata [1] ) );
BUF_X1 \AXI4Interconnect/_1935_ ( .A(\AXI4Interconnect/_0511_ ), .Z(\io_master_wdata [2] ) );
BUF_X1 \AXI4Interconnect/_1936_ ( .A(\AXI4Interconnect/_0514_ ), .Z(\io_master_wdata [3] ) );
BUF_X1 \AXI4Interconnect/_1937_ ( .A(\AXI4Interconnect/_0515_ ), .Z(\io_master_wdata [4] ) );
BUF_X1 \AXI4Interconnect/_1938_ ( .A(\AXI4Interconnect/_0516_ ), .Z(\io_master_wdata [5] ) );
BUF_X1 \AXI4Interconnect/_1939_ ( .A(\AXI4Interconnect/_0517_ ), .Z(\io_master_wdata [6] ) );
BUF_X1 \AXI4Interconnect/_1940_ ( .A(\AXI4Interconnect/_0518_ ), .Z(\io_master_wdata [7] ) );
BUF_X1 \AXI4Interconnect/_1941_ ( .A(\AXI4Interconnect/_0519_ ), .Z(\io_master_wdata [8] ) );
BUF_X1 \AXI4Interconnect/_1942_ ( .A(\AXI4Interconnect/_0520_ ), .Z(\io_master_wdata [9] ) );
BUF_X1 \AXI4Interconnect/_1943_ ( .A(\AXI4Interconnect/_0490_ ), .Z(\io_master_wdata [10] ) );
BUF_X1 \AXI4Interconnect/_1944_ ( .A(\AXI4Interconnect/_0491_ ), .Z(\io_master_wdata [11] ) );
BUF_X1 \AXI4Interconnect/_1945_ ( .A(\AXI4Interconnect/_0492_ ), .Z(\io_master_wdata [12] ) );
BUF_X1 \AXI4Interconnect/_1946_ ( .A(\AXI4Interconnect/_0493_ ), .Z(\io_master_wdata [13] ) );
BUF_X1 \AXI4Interconnect/_1947_ ( .A(\AXI4Interconnect/_0494_ ), .Z(\io_master_wdata [14] ) );
BUF_X1 \AXI4Interconnect/_1948_ ( .A(\AXI4Interconnect/_0495_ ), .Z(\io_master_wdata [15] ) );
BUF_X1 \AXI4Interconnect/_1949_ ( .A(\AXI4Interconnect/_0496_ ), .Z(\io_master_wdata [16] ) );
BUF_X1 \AXI4Interconnect/_1950_ ( .A(\AXI4Interconnect/_0497_ ), .Z(\io_master_wdata [17] ) );
BUF_X1 \AXI4Interconnect/_1951_ ( .A(\AXI4Interconnect/_0498_ ), .Z(\io_master_wdata [18] ) );
BUF_X1 \AXI4Interconnect/_1952_ ( .A(\AXI4Interconnect/_0499_ ), .Z(\io_master_wdata [19] ) );
BUF_X1 \AXI4Interconnect/_1953_ ( .A(\AXI4Interconnect/_0501_ ), .Z(\io_master_wdata [20] ) );
BUF_X1 \AXI4Interconnect/_1954_ ( .A(\AXI4Interconnect/_0502_ ), .Z(\io_master_wdata [21] ) );
BUF_X1 \AXI4Interconnect/_1955_ ( .A(\AXI4Interconnect/_0503_ ), .Z(\io_master_wdata [22] ) );
BUF_X1 \AXI4Interconnect/_1956_ ( .A(\AXI4Interconnect/_0504_ ), .Z(\io_master_wdata [23] ) );
BUF_X1 \AXI4Interconnect/_1957_ ( .A(\AXI4Interconnect/_0505_ ), .Z(\io_master_wdata [24] ) );
BUF_X1 \AXI4Interconnect/_1958_ ( .A(\AXI4Interconnect/_0506_ ), .Z(\io_master_wdata [25] ) );
BUF_X1 \AXI4Interconnect/_1959_ ( .A(\AXI4Interconnect/_0507_ ), .Z(\io_master_wdata [26] ) );
BUF_X1 \AXI4Interconnect/_1960_ ( .A(\AXI4Interconnect/_0508_ ), .Z(\io_master_wdata [27] ) );
BUF_X1 \AXI4Interconnect/_1961_ ( .A(\AXI4Interconnect/_0509_ ), .Z(\io_master_wdata [28] ) );
BUF_X1 \AXI4Interconnect/_1962_ ( .A(\AXI4Interconnect/_0510_ ), .Z(\io_master_wdata [29] ) );
BUF_X1 \AXI4Interconnect/_1963_ ( .A(\AXI4Interconnect/_0512_ ), .Z(\io_master_wdata [30] ) );
BUF_X1 \AXI4Interconnect/_1964_ ( .A(\AXI4Interconnect/_0513_ ), .Z(\io_master_wdata [31] ) );
BUF_X1 \AXI4Interconnect/_1965_ ( .A(\_LSU_io_master_wstrb [0] ), .Z(\AXI4Interconnect/_0228_ ) );
BUF_X1 \AXI4Interconnect/_1966_ ( .A(\AXI4Interconnect/_0523_ ), .Z(\io_master_wstrb [0] ) );
BUF_X1 \AXI4Interconnect/_1967_ ( .A(\_LSU_io_master_wstrb [1] ), .Z(\AXI4Interconnect/_0229_ ) );
BUF_X1 \AXI4Interconnect/_1968_ ( .A(\AXI4Interconnect/_0524_ ), .Z(\io_master_wstrb [1] ) );
BUF_X1 \AXI4Interconnect/_1969_ ( .A(\_LSU_io_master_wstrb [2] ), .Z(\AXI4Interconnect/_0230_ ) );
BUF_X1 \AXI4Interconnect/_1970_ ( .A(\AXI4Interconnect/_0525_ ), .Z(\io_master_wstrb [2] ) );
BUF_X1 \AXI4Interconnect/_1971_ ( .A(\_LSU_io_master_wstrb [3] ), .Z(\AXI4Interconnect/_0231_ ) );
BUF_X1 \AXI4Interconnect/_1972_ ( .A(\AXI4Interconnect/_0526_ ), .Z(\io_master_wstrb [3] ) );
BUF_X1 \AXI4Interconnect/_1973_ ( .A(\AXI4Interconnect/_0375_ ), .Z(\io_master_araddr [0] ) );
BUF_X1 \AXI4Interconnect/_1974_ ( .A(\AXI4Interconnect/_0386_ ), .Z(\io_master_araddr [1] ) );
BUF_X1 \AXI4Interconnect/_1975_ ( .A(\AXI4Interconnect/_0397_ ), .Z(\io_master_araddr [2] ) );
BUF_X1 \AXI4Interconnect/_1976_ ( .A(\AXI4Interconnect/_0400_ ), .Z(\io_master_araddr [3] ) );
BUF_X1 \AXI4Interconnect/_1977_ ( .A(\AXI4Interconnect/_0401_ ), .Z(\io_master_araddr [4] ) );
BUF_X1 \AXI4Interconnect/_1978_ ( .A(\AXI4Interconnect/_0402_ ), .Z(\io_master_araddr [5] ) );
BUF_X1 \AXI4Interconnect/_1979_ ( .A(\AXI4Interconnect/_0403_ ), .Z(\io_master_araddr [6] ) );
BUF_X1 \AXI4Interconnect/_1980_ ( .A(\AXI4Interconnect/_0404_ ), .Z(\io_master_araddr [7] ) );
BUF_X1 \AXI4Interconnect/_1981_ ( .A(\AXI4Interconnect/_0405_ ), .Z(\io_master_araddr [8] ) );
BUF_X1 \AXI4Interconnect/_1982_ ( .A(\AXI4Interconnect/_0406_ ), .Z(\io_master_araddr [9] ) );
BUF_X1 \AXI4Interconnect/_1983_ ( .A(\AXI4Interconnect/_0376_ ), .Z(\io_master_araddr [10] ) );
BUF_X1 \AXI4Interconnect/_1984_ ( .A(\AXI4Interconnect/_0377_ ), .Z(\io_master_araddr [11] ) );
BUF_X1 \AXI4Interconnect/_1985_ ( .A(\AXI4Interconnect/_0378_ ), .Z(\io_master_araddr [12] ) );
BUF_X1 \AXI4Interconnect/_1986_ ( .A(\AXI4Interconnect/_0379_ ), .Z(\io_master_araddr [13] ) );
BUF_X1 \AXI4Interconnect/_1987_ ( .A(\AXI4Interconnect/_0380_ ), .Z(\io_master_araddr [14] ) );
BUF_X1 \AXI4Interconnect/_1988_ ( .A(\AXI4Interconnect/_0381_ ), .Z(\io_master_araddr [15] ) );
BUF_X1 \AXI4Interconnect/_1989_ ( .A(\AXI4Interconnect/_0382_ ), .Z(\io_master_araddr [16] ) );
BUF_X1 \AXI4Interconnect/_1990_ ( .A(\AXI4Interconnect/_0383_ ), .Z(\io_master_araddr [17] ) );
BUF_X1 \AXI4Interconnect/_1991_ ( .A(\AXI4Interconnect/_0384_ ), .Z(\io_master_araddr [18] ) );
BUF_X1 \AXI4Interconnect/_1992_ ( .A(\AXI4Interconnect/_0385_ ), .Z(\io_master_araddr [19] ) );
BUF_X1 \AXI4Interconnect/_1993_ ( .A(\AXI4Interconnect/_0387_ ), .Z(\io_master_araddr [20] ) );
BUF_X1 \AXI4Interconnect/_1994_ ( .A(\AXI4Interconnect/_0388_ ), .Z(\io_master_araddr [21] ) );
BUF_X1 \AXI4Interconnect/_1995_ ( .A(\AXI4Interconnect/_0389_ ), .Z(\io_master_araddr [22] ) );
BUF_X1 \AXI4Interconnect/_1996_ ( .A(\AXI4Interconnect/_0390_ ), .Z(\io_master_araddr [23] ) );
BUF_X1 \AXI4Interconnect/_1997_ ( .A(\AXI4Interconnect/_0391_ ), .Z(\io_master_araddr [24] ) );
BUF_X1 \AXI4Interconnect/_1998_ ( .A(\AXI4Interconnect/_0392_ ), .Z(\io_master_araddr [25] ) );
BUF_X1 \AXI4Interconnect/_1999_ ( .A(\AXI4Interconnect/_0393_ ), .Z(\io_master_araddr [26] ) );
BUF_X1 \AXI4Interconnect/_2000_ ( .A(\AXI4Interconnect/_0394_ ), .Z(\io_master_araddr [27] ) );
BUF_X1 \AXI4Interconnect/_2001_ ( .A(\AXI4Interconnect/_0395_ ), .Z(\io_master_araddr [28] ) );
BUF_X1 \AXI4Interconnect/_2002_ ( .A(\AXI4Interconnect/_0396_ ), .Z(\io_master_araddr [29] ) );
BUF_X1 \AXI4Interconnect/_2003_ ( .A(\AXI4Interconnect/_0398_ ), .Z(\io_master_araddr [30] ) );
BUF_X1 \AXI4Interconnect/_2004_ ( .A(\AXI4Interconnect/_0399_ ), .Z(\io_master_araddr [31] ) );
BUF_X1 \AXI4Interconnect/_2005_ ( .A(\_LSU_io_master_awsize [0] ), .Z(\AXI4Interconnect/_0150_ ) );
BUF_X1 \AXI4Interconnect/_2006_ ( .A(\AXI4Interconnect/_0445_ ), .Z(\io_master_awsize [0] ) );
BUF_X1 \AXI4Interconnect/_2007_ ( .A(\_LSU_io_master_awsize [1] ), .Z(\AXI4Interconnect/_0151_ ) );
BUF_X1 \AXI4Interconnect/_2008_ ( .A(\AXI4Interconnect/_0446_ ), .Z(\io_master_awsize [1] ) );
BUF_X1 \AXI4Interconnect/_2009_ ( .A(\_LSU_io_master_awsize [2] ), .Z(\AXI4Interconnect/_0152_ ) );
BUF_X1 \AXI4Interconnect/_2010_ ( .A(\AXI4Interconnect/_0447_ ), .Z(\io_master_awsize [2] ) );
BUF_X1 \AXI4Interconnect/_2011_ ( .A(\_LSU_io_master_arsize [0] ), .Z(\AXI4Interconnect/_0113_ ) );
BUF_X1 \AXI4Interconnect/_2012_ ( .A(\AXI4Interconnect/_0408_ ), .Z(\io_master_arsize [0] ) );
BUF_X1 \AXI4Interconnect/_2013_ ( .A(\_LSU_io_master_arsize [1] ), .Z(\AXI4Interconnect/_0114_ ) );
BUF_X1 \AXI4Interconnect/_2014_ ( .A(\AXI4Interconnect/_0409_ ), .Z(\io_master_arsize [1] ) );
BUF_X1 \AXI4Interconnect/_2015_ ( .A(\_LSU_io_master_arsize [2] ), .Z(\AXI4Interconnect/_0115_ ) );
BUF_X1 \AXI4Interconnect/_2016_ ( .A(\AXI4Interconnect/_0410_ ), .Z(\io_master_arsize [2] ) );
BUF_X1 \AXI4Interconnect/_2017_ ( .A(_CLINT_io_rvalid ), .Z(\AXI4Interconnect/_0340_ ) );
BUF_X1 \AXI4Interconnect/_2018_ ( .A(io_master_rvalid ), .Z(\AXI4Interconnect/_0488_ ) );
BUF_X1 \AXI4Interconnect/_2019_ ( .A(_IFU_io_master_rready ), .Z(\AXI4Interconnect/_0076_ ) );
BUF_X1 \AXI4Interconnect/_2020_ ( .A(_LSU_io_master_rready ), .Z(\AXI4Interconnect/_0190_ ) );
BUF_X1 \AXI4Interconnect/_2021_ ( .A(_LSU_io_master_wvalid ), .Z(\AXI4Interconnect/_0232_ ) );
BUF_X1 \AXI4Interconnect/_2022_ ( .A(_CLINT_io_wready ), .Z(\AXI4Interconnect/_0373_ ) );
BUF_X1 \AXI4Interconnect/_2023_ ( .A(io_master_wready ), .Z(\AXI4Interconnect/_0522_ ) );
BUF_X1 \AXI4Interconnect/_2024_ ( .A(_IFU_io_master_arvalid ), .Z(\AXI4Interconnect/_0043_ ) );
BUF_X1 \AXI4Interconnect/_2025_ ( .A(_LSU_io_master_awvalid ), .Z(\AXI4Interconnect/_0153_ ) );
BUF_X1 \AXI4Interconnect/_2026_ ( .A(_LSU_io_master_arvalid ), .Z(\AXI4Interconnect/_0116_ ) );
BUF_X1 \AXI4Interconnect/_2027_ ( .A(_CLINT_io_bvalid ), .Z(\AXI4Interconnect/_0304_ ) );
BUF_X1 \AXI4Interconnect/_2028_ ( .A(io_master_bvalid ), .Z(\AXI4Interconnect/_0452_ ) );
BUF_X1 \AXI4Interconnect/_2029_ ( .A(_LSU_io_master_bready ), .Z(\AXI4Interconnect/_0154_ ) );
BUF_X1 \AXI4Interconnect/_2030_ ( .A(_CLINT_io_arready ), .Z(\AXI4Interconnect/_0265_ ) );
BUF_X1 \AXI4Interconnect/_2031_ ( .A(io_master_arready ), .Z(\AXI4Interconnect/_0407_ ) );
BUF_X1 \AXI4Interconnect/_2032_ ( .A(\AXI4Interconnect/_0042_ ), .Z(_AXI4Interconnect_io_fanIn_0_arready ) );
BUF_X1 \AXI4Interconnect/_2033_ ( .A(\AXI4Interconnect/_0079_ ), .Z(_AXI4Interconnect_io_fanIn_0_rvalid ) );
BUF_X1 \AXI4Interconnect/_2034_ ( .A(_CLINT_io_awready ), .Z(\AXI4Interconnect/_0299_ ) );
BUF_X1 \AXI4Interconnect/_2035_ ( .A(io_master_awready ), .Z(\AXI4Interconnect/_0444_ ) );
BUF_X1 \AXI4Interconnect/_2036_ ( .A(\AXI4Interconnect/_0149_ ), .Z(_AXI4Interconnect_io_fanIn_1_awready ) );
BUF_X1 \AXI4Interconnect/_2037_ ( .A(\AXI4Interconnect/_0227_ ), .Z(_AXI4Interconnect_io_fanIn_1_wready ) );
BUF_X1 \AXI4Interconnect/_2038_ ( .A(\AXI4Interconnect/_0157_ ), .Z(_AXI4Interconnect_io_fanIn_1_bvalid ) );
BUF_X1 \AXI4Interconnect/_2039_ ( .A(\AXI4Interconnect/_0112_ ), .Z(_AXI4Interconnect_io_fanIn_1_arready ) );
BUF_X1 \AXI4Interconnect/_2040_ ( .A(\AXI4Interconnect/_0193_ ), .Z(_AXI4Interconnect_io_fanIn_1_rvalid ) );
BUF_X1 \AXI4Interconnect/_2041_ ( .A(\AXI4Interconnect/_0300_ ), .Z(_AXI4Interconnect_io_fanOut_0_awvalid ) );
BUF_X1 \AXI4Interconnect/_2042_ ( .A(\AXI4Interconnect/_0374_ ), .Z(_AXI4Interconnect_io_fanOut_0_wvalid ) );
BUF_X1 \AXI4Interconnect/_2043_ ( .A(\AXI4Interconnect/_0301_ ), .Z(_AXI4Interconnect_io_fanOut_0_bready ) );
BUF_X1 \AXI4Interconnect/_2044_ ( .A(\AXI4Interconnect/_0266_ ), .Z(_AXI4Interconnect_io_fanOut_0_arvalid ) );
BUF_X1 \AXI4Interconnect/_2045_ ( .A(\AXI4Interconnect/_0337_ ), .Z(_AXI4Interconnect_io_fanOut_0_rready ) );
BUF_X1 \AXI4Interconnect/_2046_ ( .A(\AXI4Interconnect/_0448_ ), .Z(io_master_awvalid ) );
BUF_X1 \AXI4Interconnect/_2047_ ( .A(\AXI4Interconnect/_0527_ ), .Z(io_master_wvalid ) );
BUF_X1 \AXI4Interconnect/_2048_ ( .A(\AXI4Interconnect/_0449_ ), .Z(io_master_bready ) );
BUF_X1 \AXI4Interconnect/_2049_ ( .A(\AXI4Interconnect/_0411_ ), .Z(io_master_arvalid ) );
BUF_X1 \AXI4Interconnect/_2050_ ( .A(\AXI4Interconnect/_0485_ ), .Z(io_master_rready ) );
BUF_X1 \AXI4Interconnect/_2051_ ( .A(_LSU_io_master_wlast ), .Z(\AXI4Interconnect/_0226_ ) );
BUF_X1 \AXI4Interconnect/_2052_ ( .A(\AXI4Interconnect/_0521_ ), .Z(io_master_wlast ) );
BUF_X1 \AXI4Interconnect/_2053_ ( .A(reset ), .Z(\AXI4Interconnect/_0870_ ) );
BUF_X1 \AXI4Interconnect/_2054_ ( .A(\AXI4Interconnect/_0006_ ), .Z(\AXI4Interconnect/_0877_ ) );
BUF_X1 \AXI4Interconnect/_2055_ ( .A(\AXI4Interconnect/_0007_ ), .Z(\AXI4Interconnect/_0878_ ) );
BUF_X1 \AXI4Interconnect/_2056_ ( .A(\AXI4Interconnect/_0008_ ), .Z(\AXI4Interconnect/_0879_ ) );
BUF_X1 \AXI4Interconnect/_2057_ ( .A(\AXI4Interconnect/_0009_ ), .Z(\AXI4Interconnect/_0880_ ) );
NOR2_X1 \CLINT/_0838_ ( .A1(\CLINT/_0578_ ), .A2(\CLINT/_0579_ ), .ZN(\CLINT/_0237_ ) );
AND2_X1 \CLINT/_0839_ ( .A1(\CLINT/_0237_ ), .A2(\CLINT/_0580_ ), .ZN(\CLINT/_0170_ ) );
AND3_X1 \CLINT/_0840_ ( .A1(\CLINT/_0578_ ), .A2(\CLINT/_0579_ ), .A3(\CLINT/_0001_ ), .ZN(\CLINT/_0135_ ) );
OR2_X1 \CLINT/_0841_ ( .A1(\CLINT/_0569_ ), .A2(\CLINT/_0568_ ), .ZN(\CLINT/_0238_ ) );
OR3_X1 \CLINT/_0842_ ( .A1(\CLINT/_0238_ ), .A2(\CLINT/_0566_ ), .A3(\CLINT/_0565_ ), .ZN(\CLINT/_0239_ ) );
INV_X1 \CLINT/_0843_ ( .A(\CLINT/_0561_ ), .ZN(\CLINT/_0240_ ) );
NAND2_X1 \CLINT/_0844_ ( .A1(\CLINT/_0240_ ), .A2(\CLINT/_0562_ ), .ZN(\CLINT/_0241_ ) );
NOR4_X1 \CLINT/_0845_ ( .A1(\CLINT/_0239_ ), .A2(\CLINT/_0564_ ), .A3(\CLINT/_0563_ ), .A4(\CLINT/_0241_ ), .ZN(\CLINT/_0242_ ) );
NOR4_X1 \CLINT/_0846_ ( .A1(\CLINT/_0558_ ), .A2(\CLINT/_0557_ ), .A3(\CLINT/_0560_ ), .A4(\CLINT/_0559_ ), .ZN(\CLINT/_0243_ ) );
NOR4_X1 \CLINT/_0847_ ( .A1(\CLINT/_0554_ ), .A2(\CLINT/_0553_ ), .A3(\CLINT/_0556_ ), .A4(\CLINT/_0555_ ), .ZN(\CLINT/_0244_ ) );
AND2_X1 \CLINT/_0848_ ( .A1(\CLINT/_0243_ ), .A2(\CLINT/_0244_ ), .ZN(\CLINT/_0245_ ) );
AND2_X1 \CLINT/_0849_ ( .A1(\CLINT/_0242_ ), .A2(\CLINT/_0245_ ), .ZN(\CLINT/_0246_ ) );
BUF_X4 \CLINT/_0850_ ( .A(\CLINT/_0246_ ), .Z(\CLINT/_0247_ ) );
BUF_X4 \CLINT/_0851_ ( .A(\CLINT/_0247_ ), .Z(\CLINT/_0248_ ) );
OR4_X1 \CLINT/_0852_ ( .A1(\CLINT/_0550_ ), .A2(\CLINT/_0549_ ), .A3(\CLINT/_0552_ ), .A4(\CLINT/_0551_ ), .ZN(\CLINT/_0249_ ) );
NOR3_X1 \CLINT/_0853_ ( .A1(\CLINT/_0249_ ), .A2(\CLINT/_0548_ ), .A3(\CLINT/_0547_ ), .ZN(\CLINT/_0250_ ) );
BUF_X4 \CLINT/_0854_ ( .A(\CLINT/_0250_ ), .Z(\CLINT/_0251_ ) );
BUF_X4 \CLINT/_0855_ ( .A(\CLINT/_0251_ ), .Z(\CLINT/_0252_ ) );
OR4_X1 \CLINT/_0856_ ( .A1(\CLINT/_0570_ ), .A2(\CLINT/_0572_ ), .A3(\CLINT/_0571_ ), .A4(\CLINT/_0574_ ), .ZN(\CLINT/_0253_ ) );
OR3_X1 \CLINT/_0857_ ( .A1(\CLINT/_0573_ ), .A2(\CLINT/_0576_ ), .A3(\CLINT/_0575_ ), .ZN(\CLINT/_0254_ ) );
NOR2_X1 \CLINT/_0858_ ( .A1(\CLINT/_0253_ ), .A2(\CLINT/_0254_ ), .ZN(\CLINT/_0255_ ) );
AND3_X2 \CLINT/_0859_ ( .A1(\CLINT/_0255_ ), .A2(\CLINT/_0567_ ), .A3(\CLINT/_0170_ ), .ZN(\CLINT/_0256_ ) );
BUF_X4 \CLINT/_0860_ ( .A(\CLINT/_0256_ ), .Z(\CLINT/_0257_ ) );
NAND4_X1 \CLINT/_0861_ ( .A1(\CLINT/_0248_ ), .A2(\CLINT/_0198_ ), .A3(\CLINT/_0252_ ), .A4(\CLINT/_0257_ ), .ZN(\CLINT/_0258_ ) );
BUF_X4 \CLINT/_0862_ ( .A(\CLINT/_0247_ ), .Z(\CLINT/_0259_ ) );
BUF_X4 \CLINT/_0863_ ( .A(\CLINT/_0251_ ), .Z(\CLINT/_0260_ ) );
INV_X1 \CLINT/_0864_ ( .A(\CLINT/_0580_ ), .ZN(\CLINT/_0261_ ) );
OR4_X1 \CLINT/_0865_ ( .A1(\CLINT/_0578_ ), .A2(\CLINT/_0261_ ), .A3(\CLINT/_0579_ ), .A4(\CLINT/_0567_ ), .ZN(\CLINT/_0262_ ) );
NOR3_X4 \CLINT/_0866_ ( .A1(\CLINT/_0262_ ), .A2(\CLINT/_0253_ ), .A3(\CLINT/_0254_ ), .ZN(\CLINT/_0263_ ) );
BUF_X4 \CLINT/_0867_ ( .A(\CLINT/_0263_ ), .Z(\CLINT/_0264_ ) );
NAND4_X1 \CLINT/_0868_ ( .A1(\CLINT/_0259_ ), .A2(\CLINT/_0173_ ), .A3(\CLINT/_0260_ ), .A4(\CLINT/_0264_ ), .ZN(\CLINT/_0265_ ) );
NAND2_X1 \CLINT/_0869_ ( .A1(\CLINT/_0258_ ), .A2(\CLINT/_0265_ ), .ZN(\CLINT/_0136_ ) );
NAND4_X1 \CLINT/_0870_ ( .A1(\CLINT/_0248_ ), .A2(\CLINT/_0199_ ), .A3(\CLINT/_0252_ ), .A4(\CLINT/_0257_ ), .ZN(\CLINT/_0266_ ) );
NAND4_X1 \CLINT/_0871_ ( .A1(\CLINT/_0259_ ), .A2(\CLINT/_0184_ ), .A3(\CLINT/_0260_ ), .A4(\CLINT/_0264_ ), .ZN(\CLINT/_0267_ ) );
NAND2_X1 \CLINT/_0872_ ( .A1(\CLINT/_0266_ ), .A2(\CLINT/_0267_ ), .ZN(\CLINT/_0147_ ) );
NAND4_X1 \CLINT/_0873_ ( .A1(\CLINT/_0248_ ), .A2(\CLINT/_0200_ ), .A3(\CLINT/_0252_ ), .A4(\CLINT/_0257_ ), .ZN(\CLINT/_0268_ ) );
NAND4_X1 \CLINT/_0874_ ( .A1(\CLINT/_0259_ ), .A2(\CLINT/_0195_ ), .A3(\CLINT/_0260_ ), .A4(\CLINT/_0264_ ), .ZN(\CLINT/_0269_ ) );
NAND2_X1 \CLINT/_0875_ ( .A1(\CLINT/_0268_ ), .A2(\CLINT/_0269_ ), .ZN(\CLINT/_0158_ ) );
NAND4_X1 \CLINT/_0876_ ( .A1(\CLINT/_0248_ ), .A2(\CLINT/_0201_ ), .A3(\CLINT/_0252_ ), .A4(\CLINT/_0257_ ), .ZN(\CLINT/_0270_ ) );
NAND4_X1 \CLINT/_0877_ ( .A1(\CLINT/_0259_ ), .A2(\CLINT/_0206_ ), .A3(\CLINT/_0260_ ), .A4(\CLINT/_0264_ ), .ZN(\CLINT/_0271_ ) );
NAND2_X1 \CLINT/_0878_ ( .A1(\CLINT/_0270_ ), .A2(\CLINT/_0271_ ), .ZN(\CLINT/_0161_ ) );
NAND4_X1 \CLINT/_0879_ ( .A1(\CLINT/_0248_ ), .A2(\CLINT/_0202_ ), .A3(\CLINT/_0252_ ), .A4(\CLINT/_0257_ ), .ZN(\CLINT/_0272_ ) );
NAND4_X1 \CLINT/_0880_ ( .A1(\CLINT/_0259_ ), .A2(\CLINT/_0217_ ), .A3(\CLINT/_0260_ ), .A4(\CLINT/_0264_ ), .ZN(\CLINT/_0273_ ) );
NAND2_X1 \CLINT/_0881_ ( .A1(\CLINT/_0272_ ), .A2(\CLINT/_0273_ ), .ZN(\CLINT/_0162_ ) );
NAND4_X1 \CLINT/_0882_ ( .A1(\CLINT/_0248_ ), .A2(\CLINT/_0203_ ), .A3(\CLINT/_0252_ ), .A4(\CLINT/_0257_ ), .ZN(\CLINT/_0274_ ) );
NAND4_X1 \CLINT/_0883_ ( .A1(\CLINT/_0259_ ), .A2(\CLINT/_0228_ ), .A3(\CLINT/_0260_ ), .A4(\CLINT/_0264_ ), .ZN(\CLINT/_0275_ ) );
NAND2_X1 \CLINT/_0884_ ( .A1(\CLINT/_0274_ ), .A2(\CLINT/_0275_ ), .ZN(\CLINT/_0163_ ) );
NAND4_X1 \CLINT/_0885_ ( .A1(\CLINT/_0248_ ), .A2(\CLINT/_0204_ ), .A3(\CLINT/_0252_ ), .A4(\CLINT/_0257_ ), .ZN(\CLINT/_0276_ ) );
NAND4_X1 \CLINT/_0886_ ( .A1(\CLINT/_0259_ ), .A2(\CLINT/_0233_ ), .A3(\CLINT/_0260_ ), .A4(\CLINT/_0264_ ), .ZN(\CLINT/_0277_ ) );
NAND2_X1 \CLINT/_0887_ ( .A1(\CLINT/_0276_ ), .A2(\CLINT/_0277_ ), .ZN(\CLINT/_0164_ ) );
NAND4_X1 \CLINT/_0888_ ( .A1(\CLINT/_0248_ ), .A2(\CLINT/_0205_ ), .A3(\CLINT/_0252_ ), .A4(\CLINT/_0257_ ), .ZN(\CLINT/_0278_ ) );
NAND4_X1 \CLINT/_0889_ ( .A1(\CLINT/_0259_ ), .A2(\CLINT/_0234_ ), .A3(\CLINT/_0260_ ), .A4(\CLINT/_0264_ ), .ZN(\CLINT/_0279_ ) );
NAND2_X1 \CLINT/_0890_ ( .A1(\CLINT/_0278_ ), .A2(\CLINT/_0279_ ), .ZN(\CLINT/_0165_ ) );
NAND4_X1 \CLINT/_0891_ ( .A1(\CLINT/_0248_ ), .A2(\CLINT/_0207_ ), .A3(\CLINT/_0252_ ), .A4(\CLINT/_0257_ ), .ZN(\CLINT/_0280_ ) );
BUF_X4 \CLINT/_0892_ ( .A(\CLINT/_0247_ ), .Z(\CLINT/_0281_ ) );
BUF_X4 \CLINT/_0893_ ( .A(\CLINT/_0251_ ), .Z(\CLINT/_0282_ ) );
NAND4_X1 \CLINT/_0894_ ( .A1(\CLINT/_0281_ ), .A2(\CLINT/_0235_ ), .A3(\CLINT/_0282_ ), .A4(\CLINT/_0264_ ), .ZN(\CLINT/_0283_ ) );
NAND2_X1 \CLINT/_0895_ ( .A1(\CLINT/_0280_ ), .A2(\CLINT/_0283_ ), .ZN(\CLINT/_0166_ ) );
NAND4_X1 \CLINT/_0896_ ( .A1(\CLINT/_0248_ ), .A2(\CLINT/_0208_ ), .A3(\CLINT/_0252_ ), .A4(\CLINT/_0257_ ), .ZN(\CLINT/_0284_ ) );
NAND4_X1 \CLINT/_0897_ ( .A1(\CLINT/_0281_ ), .A2(\CLINT/_0236_ ), .A3(\CLINT/_0282_ ), .A4(\CLINT/_0264_ ), .ZN(\CLINT/_0285_ ) );
NAND2_X1 \CLINT/_0898_ ( .A1(\CLINT/_0284_ ), .A2(\CLINT/_0285_ ), .ZN(\CLINT/_0167_ ) );
BUF_X4 \CLINT/_0899_ ( .A(\CLINT/_0247_ ), .Z(\CLINT/_0286_ ) );
BUF_X4 \CLINT/_0900_ ( .A(\CLINT/_0251_ ), .Z(\CLINT/_0287_ ) );
BUF_X4 \CLINT/_0901_ ( .A(\CLINT/_0256_ ), .Z(\CLINT/_0288_ ) );
NAND4_X1 \CLINT/_0902_ ( .A1(\CLINT/_0286_ ), .A2(\CLINT/_0209_ ), .A3(\CLINT/_0287_ ), .A4(\CLINT/_0288_ ), .ZN(\CLINT/_0289_ ) );
BUF_X4 \CLINT/_0903_ ( .A(\CLINT/_0263_ ), .Z(\CLINT/_0290_ ) );
NAND4_X1 \CLINT/_0904_ ( .A1(\CLINT/_0281_ ), .A2(\CLINT/_0174_ ), .A3(\CLINT/_0282_ ), .A4(\CLINT/_0290_ ), .ZN(\CLINT/_0291_ ) );
NAND2_X1 \CLINT/_0905_ ( .A1(\CLINT/_0289_ ), .A2(\CLINT/_0291_ ), .ZN(\CLINT/_0137_ ) );
NAND4_X1 \CLINT/_0906_ ( .A1(\CLINT/_0286_ ), .A2(\CLINT/_0210_ ), .A3(\CLINT/_0287_ ), .A4(\CLINT/_0288_ ), .ZN(\CLINT/_0292_ ) );
NAND4_X1 \CLINT/_0907_ ( .A1(\CLINT/_0281_ ), .A2(\CLINT/_0175_ ), .A3(\CLINT/_0282_ ), .A4(\CLINT/_0290_ ), .ZN(\CLINT/_0293_ ) );
NAND2_X1 \CLINT/_0908_ ( .A1(\CLINT/_0292_ ), .A2(\CLINT/_0293_ ), .ZN(\CLINT/_0138_ ) );
NAND4_X1 \CLINT/_0909_ ( .A1(\CLINT/_0286_ ), .A2(\CLINT/_0211_ ), .A3(\CLINT/_0287_ ), .A4(\CLINT/_0288_ ), .ZN(\CLINT/_0294_ ) );
NAND4_X1 \CLINT/_0910_ ( .A1(\CLINT/_0281_ ), .A2(\CLINT/_0176_ ), .A3(\CLINT/_0282_ ), .A4(\CLINT/_0290_ ), .ZN(\CLINT/_0295_ ) );
NAND2_X1 \CLINT/_0911_ ( .A1(\CLINT/_0294_ ), .A2(\CLINT/_0295_ ), .ZN(\CLINT/_0139_ ) );
NAND4_X1 \CLINT/_0912_ ( .A1(\CLINT/_0286_ ), .A2(\CLINT/_0212_ ), .A3(\CLINT/_0287_ ), .A4(\CLINT/_0288_ ), .ZN(\CLINT/_0296_ ) );
NAND4_X1 \CLINT/_0913_ ( .A1(\CLINT/_0281_ ), .A2(\CLINT/_0177_ ), .A3(\CLINT/_0282_ ), .A4(\CLINT/_0290_ ), .ZN(\CLINT/_0297_ ) );
NAND2_X1 \CLINT/_0914_ ( .A1(\CLINT/_0296_ ), .A2(\CLINT/_0297_ ), .ZN(\CLINT/_0140_ ) );
NAND4_X1 \CLINT/_0915_ ( .A1(\CLINT/_0286_ ), .A2(\CLINT/_0213_ ), .A3(\CLINT/_0287_ ), .A4(\CLINT/_0288_ ), .ZN(\CLINT/_0298_ ) );
NAND4_X1 \CLINT/_0916_ ( .A1(\CLINT/_0281_ ), .A2(\CLINT/_0178_ ), .A3(\CLINT/_0282_ ), .A4(\CLINT/_0290_ ), .ZN(\CLINT/_0299_ ) );
NAND2_X1 \CLINT/_0917_ ( .A1(\CLINT/_0298_ ), .A2(\CLINT/_0299_ ), .ZN(\CLINT/_0141_ ) );
NAND4_X1 \CLINT/_0918_ ( .A1(\CLINT/_0286_ ), .A2(\CLINT/_0214_ ), .A3(\CLINT/_0287_ ), .A4(\CLINT/_0288_ ), .ZN(\CLINT/_0300_ ) );
NAND4_X1 \CLINT/_0919_ ( .A1(\CLINT/_0281_ ), .A2(\CLINT/_0179_ ), .A3(\CLINT/_0282_ ), .A4(\CLINT/_0290_ ), .ZN(\CLINT/_0301_ ) );
NAND2_X1 \CLINT/_0920_ ( .A1(\CLINT/_0300_ ), .A2(\CLINT/_0301_ ), .ZN(\CLINT/_0142_ ) );
NAND4_X1 \CLINT/_0921_ ( .A1(\CLINT/_0286_ ), .A2(\CLINT/_0215_ ), .A3(\CLINT/_0287_ ), .A4(\CLINT/_0288_ ), .ZN(\CLINT/_0302_ ) );
NAND4_X1 \CLINT/_0922_ ( .A1(\CLINT/_0281_ ), .A2(\CLINT/_0180_ ), .A3(\CLINT/_0282_ ), .A4(\CLINT/_0290_ ), .ZN(\CLINT/_0303_ ) );
NAND2_X1 \CLINT/_0923_ ( .A1(\CLINT/_0302_ ), .A2(\CLINT/_0303_ ), .ZN(\CLINT/_0143_ ) );
NAND4_X1 \CLINT/_0924_ ( .A1(\CLINT/_0286_ ), .A2(\CLINT/_0216_ ), .A3(\CLINT/_0287_ ), .A4(\CLINT/_0288_ ), .ZN(\CLINT/_0304_ ) );
NAND4_X1 \CLINT/_0925_ ( .A1(\CLINT/_0281_ ), .A2(\CLINT/_0181_ ), .A3(\CLINT/_0282_ ), .A4(\CLINT/_0290_ ), .ZN(\CLINT/_0305_ ) );
NAND2_X1 \CLINT/_0926_ ( .A1(\CLINT/_0304_ ), .A2(\CLINT/_0305_ ), .ZN(\CLINT/_0144_ ) );
NAND4_X1 \CLINT/_0927_ ( .A1(\CLINT/_0286_ ), .A2(\CLINT/_0218_ ), .A3(\CLINT/_0287_ ), .A4(\CLINT/_0288_ ), .ZN(\CLINT/_0306_ ) );
BUF_X4 \CLINT/_0928_ ( .A(\CLINT/_0247_ ), .Z(\CLINT/_0307_ ) );
BUF_X4 \CLINT/_0929_ ( .A(\CLINT/_0250_ ), .Z(\CLINT/_0308_ ) );
NAND4_X1 \CLINT/_0930_ ( .A1(\CLINT/_0307_ ), .A2(\CLINT/_0182_ ), .A3(\CLINT/_0308_ ), .A4(\CLINT/_0290_ ), .ZN(\CLINT/_0309_ ) );
NAND2_X1 \CLINT/_0931_ ( .A1(\CLINT/_0306_ ), .A2(\CLINT/_0309_ ), .ZN(\CLINT/_0145_ ) );
NAND4_X1 \CLINT/_0932_ ( .A1(\CLINT/_0286_ ), .A2(\CLINT/_0219_ ), .A3(\CLINT/_0287_ ), .A4(\CLINT/_0288_ ), .ZN(\CLINT/_0310_ ) );
NAND4_X1 \CLINT/_0933_ ( .A1(\CLINT/_0307_ ), .A2(\CLINT/_0183_ ), .A3(\CLINT/_0308_ ), .A4(\CLINT/_0290_ ), .ZN(\CLINT/_0311_ ) );
NAND2_X1 \CLINT/_0934_ ( .A1(\CLINT/_0310_ ), .A2(\CLINT/_0311_ ), .ZN(\CLINT/_0146_ ) );
BUF_X4 \CLINT/_0935_ ( .A(\CLINT/_0247_ ), .Z(\CLINT/_0312_ ) );
BUF_X4 \CLINT/_0936_ ( .A(\CLINT/_0251_ ), .Z(\CLINT/_0313_ ) );
BUF_X4 \CLINT/_0937_ ( .A(\CLINT/_0256_ ), .Z(\CLINT/_0314_ ) );
NAND4_X1 \CLINT/_0938_ ( .A1(\CLINT/_0312_ ), .A2(\CLINT/_0220_ ), .A3(\CLINT/_0313_ ), .A4(\CLINT/_0314_ ), .ZN(\CLINT/_0315_ ) );
BUF_X4 \CLINT/_0939_ ( .A(\CLINT/_0263_ ), .Z(\CLINT/_0316_ ) );
NAND4_X1 \CLINT/_0940_ ( .A1(\CLINT/_0307_ ), .A2(\CLINT/_0185_ ), .A3(\CLINT/_0308_ ), .A4(\CLINT/_0316_ ), .ZN(\CLINT/_0317_ ) );
NAND2_X1 \CLINT/_0941_ ( .A1(\CLINT/_0315_ ), .A2(\CLINT/_0317_ ), .ZN(\CLINT/_0148_ ) );
NAND4_X1 \CLINT/_0942_ ( .A1(\CLINT/_0312_ ), .A2(\CLINT/_0221_ ), .A3(\CLINT/_0313_ ), .A4(\CLINT/_0314_ ), .ZN(\CLINT/_0318_ ) );
NAND4_X1 \CLINT/_0943_ ( .A1(\CLINT/_0307_ ), .A2(\CLINT/_0186_ ), .A3(\CLINT/_0308_ ), .A4(\CLINT/_0316_ ), .ZN(\CLINT/_0319_ ) );
NAND2_X1 \CLINT/_0944_ ( .A1(\CLINT/_0318_ ), .A2(\CLINT/_0319_ ), .ZN(\CLINT/_0149_ ) );
NAND4_X1 \CLINT/_0945_ ( .A1(\CLINT/_0312_ ), .A2(\CLINT/_0222_ ), .A3(\CLINT/_0313_ ), .A4(\CLINT/_0314_ ), .ZN(\CLINT/_0320_ ) );
NAND4_X1 \CLINT/_0946_ ( .A1(\CLINT/_0307_ ), .A2(\CLINT/_0187_ ), .A3(\CLINT/_0308_ ), .A4(\CLINT/_0316_ ), .ZN(\CLINT/_0321_ ) );
NAND2_X1 \CLINT/_0947_ ( .A1(\CLINT/_0320_ ), .A2(\CLINT/_0321_ ), .ZN(\CLINT/_0150_ ) );
NAND4_X1 \CLINT/_0948_ ( .A1(\CLINT/_0312_ ), .A2(\CLINT/_0223_ ), .A3(\CLINT/_0313_ ), .A4(\CLINT/_0314_ ), .ZN(\CLINT/_0322_ ) );
NAND4_X1 \CLINT/_0949_ ( .A1(\CLINT/_0307_ ), .A2(\CLINT/_0188_ ), .A3(\CLINT/_0308_ ), .A4(\CLINT/_0316_ ), .ZN(\CLINT/_0323_ ) );
NAND2_X1 \CLINT/_0950_ ( .A1(\CLINT/_0322_ ), .A2(\CLINT/_0323_ ), .ZN(\CLINT/_0151_ ) );
NAND4_X1 \CLINT/_0951_ ( .A1(\CLINT/_0312_ ), .A2(\CLINT/_0224_ ), .A3(\CLINT/_0313_ ), .A4(\CLINT/_0314_ ), .ZN(\CLINT/_0324_ ) );
NAND4_X1 \CLINT/_0952_ ( .A1(\CLINT/_0307_ ), .A2(\CLINT/_0189_ ), .A3(\CLINT/_0308_ ), .A4(\CLINT/_0316_ ), .ZN(\CLINT/_0325_ ) );
NAND2_X1 \CLINT/_0953_ ( .A1(\CLINT/_0324_ ), .A2(\CLINT/_0325_ ), .ZN(\CLINT/_0152_ ) );
NAND4_X1 \CLINT/_0954_ ( .A1(\CLINT/_0312_ ), .A2(\CLINT/_0225_ ), .A3(\CLINT/_0313_ ), .A4(\CLINT/_0314_ ), .ZN(\CLINT/_0326_ ) );
NAND4_X1 \CLINT/_0955_ ( .A1(\CLINT/_0307_ ), .A2(\CLINT/_0190_ ), .A3(\CLINT/_0308_ ), .A4(\CLINT/_0316_ ), .ZN(\CLINT/_0327_ ) );
NAND2_X1 \CLINT/_0956_ ( .A1(\CLINT/_0326_ ), .A2(\CLINT/_0327_ ), .ZN(\CLINT/_0153_ ) );
NAND4_X1 \CLINT/_0957_ ( .A1(\CLINT/_0312_ ), .A2(\CLINT/_0226_ ), .A3(\CLINT/_0313_ ), .A4(\CLINT/_0314_ ), .ZN(\CLINT/_0328_ ) );
NAND4_X1 \CLINT/_0958_ ( .A1(\CLINT/_0307_ ), .A2(\CLINT/_0191_ ), .A3(\CLINT/_0308_ ), .A4(\CLINT/_0316_ ), .ZN(\CLINT/_0329_ ) );
NAND2_X1 \CLINT/_0959_ ( .A1(\CLINT/_0328_ ), .A2(\CLINT/_0329_ ), .ZN(\CLINT/_0154_ ) );
NAND4_X1 \CLINT/_0960_ ( .A1(\CLINT/_0312_ ), .A2(\CLINT/_0227_ ), .A3(\CLINT/_0313_ ), .A4(\CLINT/_0314_ ), .ZN(\CLINT/_0330_ ) );
NAND4_X1 \CLINT/_0961_ ( .A1(\CLINT/_0307_ ), .A2(\CLINT/_0192_ ), .A3(\CLINT/_0308_ ), .A4(\CLINT/_0316_ ), .ZN(\CLINT/_0331_ ) );
NAND2_X1 \CLINT/_0962_ ( .A1(\CLINT/_0330_ ), .A2(\CLINT/_0331_ ), .ZN(\CLINT/_0155_ ) );
NAND4_X1 \CLINT/_0963_ ( .A1(\CLINT/_0312_ ), .A2(\CLINT/_0229_ ), .A3(\CLINT/_0313_ ), .A4(\CLINT/_0314_ ), .ZN(\CLINT/_0332_ ) );
NAND4_X1 \CLINT/_0964_ ( .A1(\CLINT/_0247_ ), .A2(\CLINT/_0193_ ), .A3(\CLINT/_0251_ ), .A4(\CLINT/_0316_ ), .ZN(\CLINT/_0333_ ) );
NAND2_X1 \CLINT/_0965_ ( .A1(\CLINT/_0332_ ), .A2(\CLINT/_0333_ ), .ZN(\CLINT/_0156_ ) );
NAND4_X1 \CLINT/_0966_ ( .A1(\CLINT/_0312_ ), .A2(\CLINT/_0230_ ), .A3(\CLINT/_0313_ ), .A4(\CLINT/_0314_ ), .ZN(\CLINT/_0334_ ) );
NAND4_X1 \CLINT/_0967_ ( .A1(\CLINT/_0247_ ), .A2(\CLINT/_0194_ ), .A3(\CLINT/_0251_ ), .A4(\CLINT/_0316_ ), .ZN(\CLINT/_0335_ ) );
NAND2_X1 \CLINT/_0968_ ( .A1(\CLINT/_0334_ ), .A2(\CLINT/_0335_ ), .ZN(\CLINT/_0157_ ) );
NAND4_X1 \CLINT/_0969_ ( .A1(\CLINT/_0259_ ), .A2(\CLINT/_0231_ ), .A3(\CLINT/_0260_ ), .A4(\CLINT/_0256_ ), .ZN(\CLINT/_0336_ ) );
NAND4_X1 \CLINT/_0970_ ( .A1(\CLINT/_0247_ ), .A2(\CLINT/_0196_ ), .A3(\CLINT/_0251_ ), .A4(\CLINT/_0263_ ), .ZN(\CLINT/_0337_ ) );
NAND2_X1 \CLINT/_0971_ ( .A1(\CLINT/_0336_ ), .A2(\CLINT/_0337_ ), .ZN(\CLINT/_0159_ ) );
NAND4_X1 \CLINT/_0972_ ( .A1(\CLINT/_0259_ ), .A2(\CLINT/_0232_ ), .A3(\CLINT/_0260_ ), .A4(\CLINT/_0256_ ), .ZN(\CLINT/_0338_ ) );
NAND4_X1 \CLINT/_0973_ ( .A1(\CLINT/_0247_ ), .A2(\CLINT/_0197_ ), .A3(\CLINT/_0251_ ), .A4(\CLINT/_0263_ ), .ZN(\CLINT/_0339_ ) );
NAND2_X1 \CLINT/_0974_ ( .A1(\CLINT/_0338_ ), .A2(\CLINT/_0339_ ), .ZN(\CLINT/_0160_ ) );
AND2_X1 \CLINT/_0975_ ( .A1(\CLINT/_0237_ ), .A2(\CLINT/_0261_ ), .ZN(\CLINT/_0130_ ) );
AND2_X1 \CLINT/_0976_ ( .A1(\CLINT/_0578_ ), .A2(\CLINT/_0001_ ), .ZN(\CLINT/_0340_ ) );
INV_X1 \CLINT/_0977_ ( .A(\CLINT/_0579_ ), .ZN(\CLINT/_0341_ ) );
AND2_X1 \CLINT/_0978_ ( .A1(\CLINT/_0340_ ), .A2(\CLINT/_0341_ ), .ZN(\CLINT/_0342_ ) );
OR2_X1 \CLINT/_0979_ ( .A1(\CLINT/_0342_ ), .A2(\CLINT/_0130_ ), .ZN(\CLINT/_0132_ ) );
NAND2_X1 \CLINT/_0980_ ( .A1(\CLINT/_0579_ ), .A2(\CLINT/_0001_ ), .ZN(\CLINT/_0343_ ) );
NOR2_X1 \CLINT/_0981_ ( .A1(\CLINT/_0343_ ), .A2(\CLINT/_0578_ ), .ZN(\CLINT/_0344_ ) );
OR2_X1 \CLINT/_0982_ ( .A1(\CLINT/_0130_ ), .A2(\CLINT/_0344_ ), .ZN(\CLINT/_0171_ ) );
NAND4_X1 \CLINT/_0983_ ( .A1(\CLINT/_0242_ ), .A2(\CLINT/_0251_ ), .A3(\CLINT/_0245_ ), .A4(\CLINT/_0255_ ), .ZN(\CLINT/_0345_ ) );
AND2_X1 \CLINT/_0984_ ( .A1(\CLINT/_0345_ ), .A2(\CLINT/_0170_ ), .ZN(\CLINT/_0169_ ) );
AND2_X2 \CLINT/_0985_ ( .A1(\CLINT/_0130_ ), .A2(\CLINT/_0131_ ), .ZN(\CLINT/_0346_ ) );
BUF_X4 \CLINT/_0986_ ( .A(\CLINT/_0346_ ), .Z(\CLINT/_0347_ ) );
MUX2_X1 \CLINT/_0987_ ( .A(\CLINT/_0567_ ), .B(\CLINT/_0120_ ), .S(\CLINT/_0347_ ), .Z(\CLINT/_0005_ ) );
MUX2_X1 \CLINT/_0988_ ( .A(\CLINT/_0570_ ), .B(\CLINT/_0123_ ), .S(\CLINT/_0347_ ), .Z(\CLINT/_0006_ ) );
MUX2_X1 \CLINT/_0989_ ( .A(\CLINT/_0571_ ), .B(\CLINT/_0124_ ), .S(\CLINT/_0347_ ), .Z(\CLINT/_0007_ ) );
MUX2_X1 \CLINT/_0990_ ( .A(\CLINT/_0572_ ), .B(\CLINT/_0125_ ), .S(\CLINT/_0347_ ), .Z(\CLINT/_0008_ ) );
MUX2_X1 \CLINT/_0991_ ( .A(\CLINT/_0573_ ), .B(\CLINT/_0126_ ), .S(\CLINT/_0347_ ), .Z(\CLINT/_0009_ ) );
MUX2_X1 \CLINT/_0992_ ( .A(\CLINT/_0574_ ), .B(\CLINT/_0127_ ), .S(\CLINT/_0347_ ), .Z(\CLINT/_0010_ ) );
MUX2_X1 \CLINT/_0993_ ( .A(\CLINT/_0575_ ), .B(\CLINT/_0128_ ), .S(\CLINT/_0347_ ), .Z(\CLINT/_0011_ ) );
MUX2_X1 \CLINT/_0994_ ( .A(\CLINT/_0576_ ), .B(\CLINT/_0129_ ), .S(\CLINT/_0347_ ), .Z(\CLINT/_0012_ ) );
MUX2_X1 \CLINT/_0995_ ( .A(\CLINT/_0547_ ), .B(\CLINT/_0100_ ), .S(\CLINT/_0347_ ), .Z(\CLINT/_0013_ ) );
MUX2_X1 \CLINT/_0996_ ( .A(\CLINT/_0548_ ), .B(\CLINT/_0101_ ), .S(\CLINT/_0347_ ), .Z(\CLINT/_0014_ ) );
BUF_X4 \CLINT/_0997_ ( .A(\CLINT/_0346_ ), .Z(\CLINT/_0348_ ) );
MUX2_X1 \CLINT/_0998_ ( .A(\CLINT/_0549_ ), .B(\CLINT/_0102_ ), .S(\CLINT/_0348_ ), .Z(\CLINT/_0015_ ) );
MUX2_X1 \CLINT/_0999_ ( .A(\CLINT/_0550_ ), .B(\CLINT/_0103_ ), .S(\CLINT/_0348_ ), .Z(\CLINT/_0016_ ) );
MUX2_X1 \CLINT/_1000_ ( .A(\CLINT/_0551_ ), .B(\CLINT/_0104_ ), .S(\CLINT/_0348_ ), .Z(\CLINT/_0017_ ) );
MUX2_X1 \CLINT/_1001_ ( .A(\CLINT/_0552_ ), .B(\CLINT/_0105_ ), .S(\CLINT/_0348_ ), .Z(\CLINT/_0018_ ) );
MUX2_X1 \CLINT/_1002_ ( .A(\CLINT/_0553_ ), .B(\CLINT/_0106_ ), .S(\CLINT/_0348_ ), .Z(\CLINT/_0019_ ) );
MUX2_X1 \CLINT/_1003_ ( .A(\CLINT/_0554_ ), .B(\CLINT/_0107_ ), .S(\CLINT/_0348_ ), .Z(\CLINT/_0020_ ) );
MUX2_X1 \CLINT/_1004_ ( .A(\CLINT/_0555_ ), .B(\CLINT/_0108_ ), .S(\CLINT/_0348_ ), .Z(\CLINT/_0021_ ) );
MUX2_X1 \CLINT/_1005_ ( .A(\CLINT/_0556_ ), .B(\CLINT/_0109_ ), .S(\CLINT/_0348_ ), .Z(\CLINT/_0022_ ) );
MUX2_X1 \CLINT/_1006_ ( .A(\CLINT/_0557_ ), .B(\CLINT/_0110_ ), .S(\CLINT/_0348_ ), .Z(\CLINT/_0023_ ) );
MUX2_X1 \CLINT/_1007_ ( .A(\CLINT/_0558_ ), .B(\CLINT/_0111_ ), .S(\CLINT/_0348_ ), .Z(\CLINT/_0024_ ) );
BUF_X4 \CLINT/_1008_ ( .A(\CLINT/_0346_ ), .Z(\CLINT/_0349_ ) );
MUX2_X1 \CLINT/_1009_ ( .A(\CLINT/_0559_ ), .B(\CLINT/_0112_ ), .S(\CLINT/_0349_ ), .Z(\CLINT/_0025_ ) );
MUX2_X1 \CLINT/_1010_ ( .A(\CLINT/_0560_ ), .B(\CLINT/_0113_ ), .S(\CLINT/_0349_ ), .Z(\CLINT/_0026_ ) );
MUX2_X1 \CLINT/_1011_ ( .A(\CLINT/_0561_ ), .B(\CLINT/_0114_ ), .S(\CLINT/_0349_ ), .Z(\CLINT/_0027_ ) );
MUX2_X1 \CLINT/_1012_ ( .A(\CLINT/_0562_ ), .B(\CLINT/_0115_ ), .S(\CLINT/_0349_ ), .Z(\CLINT/_0028_ ) );
MUX2_X1 \CLINT/_1013_ ( .A(\CLINT/_0563_ ), .B(\CLINT/_0116_ ), .S(\CLINT/_0349_ ), .Z(\CLINT/_0029_ ) );
MUX2_X1 \CLINT/_1014_ ( .A(\CLINT/_0564_ ), .B(\CLINT/_0117_ ), .S(\CLINT/_0349_ ), .Z(\CLINT/_0030_ ) );
MUX2_X1 \CLINT/_1015_ ( .A(\CLINT/_0565_ ), .B(\CLINT/_0118_ ), .S(\CLINT/_0349_ ), .Z(\CLINT/_0031_ ) );
MUX2_X1 \CLINT/_1016_ ( .A(\CLINT/_0566_ ), .B(\CLINT/_0119_ ), .S(\CLINT/_0349_ ), .Z(\CLINT/_0032_ ) );
MUX2_X1 \CLINT/_1017_ ( .A(\CLINT/_0568_ ), .B(\CLINT/_0121_ ), .S(\CLINT/_0349_ ), .Z(\CLINT/_0033_ ) );
MUX2_X1 \CLINT/_1018_ ( .A(\CLINT/_0569_ ), .B(\CLINT/_0122_ ), .S(\CLINT/_0349_ ), .Z(\CLINT/_0034_ ) );
OR2_X1 \CLINT/_1019_ ( .A1(\CLINT/_0170_ ), .A2(fanout_net_7 ), .ZN(\CLINT/_0350_ ) );
INV_X1 \CLINT/_1020_ ( .A(\CLINT/_0346_ ), .ZN(\CLINT/_0351_ ) );
NAND3_X1 \CLINT/_1021_ ( .A1(\CLINT/_0351_ ), .A2(\CLINT/_0172_ ), .A3(\CLINT/_0171_ ), .ZN(\CLINT/_0352_ ) );
INV_X1 \CLINT/_1022_ ( .A(\CLINT/_0134_ ), .ZN(\CLINT/_0353_ ) );
OAI211_X2 \CLINT/_1023_ ( .A(\CLINT/_0578_ ), .B(\CLINT/_0001_ ), .C1(\CLINT/_0341_ ), .C2(\CLINT/_0353_ ), .ZN(\CLINT/_0354_ ) );
AOI21_X1 \CLINT/_1024_ ( .A(\CLINT/_0350_ ), .B1(\CLINT/_0352_ ), .B2(\CLINT/_0354_ ), .ZN(\CLINT/_0003_ ) );
NAND3_X1 \CLINT/_1025_ ( .A1(\CLINT/_0351_ ), .A2(\CLINT/_0133_ ), .A3(\CLINT/_0132_ ), .ZN(\CLINT/_0355_ ) );
AOI21_X1 \CLINT/_1026_ ( .A(\CLINT/_0344_ ), .B1(\CLINT/_0353_ ), .B2(\CLINT/_0135_ ), .ZN(\CLINT/_0356_ ) );
AOI21_X1 \CLINT/_1027_ ( .A(\CLINT/_0350_ ), .B1(\CLINT/_0355_ ), .B2(\CLINT/_0356_ ), .ZN(\CLINT/_0004_ ) );
OR4_X1 \CLINT/_1028_ ( .A1(\CLINT/_0578_ ), .A2(\CLINT/_0261_ ), .A3(\CLINT/_0579_ ), .A4(\CLINT/_0168_ ), .ZN(\CLINT/_0357_ ) );
AOI21_X1 \CLINT/_1029_ ( .A(fanout_net_7 ), .B1(\CLINT/_0351_ ), .B2(\CLINT/_0357_ ), .ZN(\CLINT/_0035_ ) );
INV_X1 \CLINT/_1030_ ( .A(fanout_net_7 ), .ZN(\CLINT/_0358_ ) );
BUF_X2 \CLINT/_1031_ ( .A(\CLINT/_0358_ ), .Z(\CLINT/_0359_ ) );
AND2_X1 \CLINT/_1032_ ( .A1(\CLINT/_0359_ ), .A2(\CLINT/_0002_ ), .ZN(\CLINT/_0036_ ) );
AND2_X4 \CLINT/_1033_ ( .A1(\CLINT/_0173_ ), .A2(\CLINT/_0184_ ), .ZN(\CLINT/_0360_ ) );
NOR2_X1 \CLINT/_1034_ ( .A1(\CLINT/_0173_ ), .A2(\CLINT/_0184_ ), .ZN(\CLINT/_0361_ ) );
NOR3_X1 \CLINT/_1035_ ( .A1(\CLINT/_0360_ ), .A2(\CLINT/_0361_ ), .A3(fanout_net_7 ), .ZN(\CLINT/_0037_ ) );
AND2_X1 \CLINT/_1036_ ( .A1(\CLINT/_0360_ ), .A2(\CLINT/_0195_ ), .ZN(\CLINT/_0362_ ) );
BUF_X4 \CLINT/_1037_ ( .A(\CLINT/_0358_ ), .Z(\CLINT/_0363_ ) );
OAI21_X1 \CLINT/_1038_ ( .A(\CLINT/_0363_ ), .B1(\CLINT/_0360_ ), .B2(\CLINT/_0195_ ), .ZN(\CLINT/_0364_ ) );
NOR2_X1 \CLINT/_1039_ ( .A1(\CLINT/_0362_ ), .A2(\CLINT/_0364_ ), .ZN(\CLINT/_0038_ ) );
AND2_X1 \CLINT/_1040_ ( .A1(\CLINT/_0362_ ), .A2(\CLINT/_0206_ ), .ZN(\CLINT/_0365_ ) );
AOI21_X1 \CLINT/_1041_ ( .A(\CLINT/_0206_ ), .B1(\CLINT/_0360_ ), .B2(\CLINT/_0195_ ), .ZN(\CLINT/_0366_ ) );
NOR3_X1 \CLINT/_1042_ ( .A1(\CLINT/_0365_ ), .A2(fanout_net_7 ), .A3(\CLINT/_0366_ ), .ZN(\CLINT/_0039_ ) );
OAI21_X1 \CLINT/_1043_ ( .A(\CLINT/_0358_ ), .B1(\CLINT/_0365_ ), .B2(\CLINT/_0217_ ), .ZN(\CLINT/_0367_ ) );
AOI21_X1 \CLINT/_1044_ ( .A(\CLINT/_0367_ ), .B1(\CLINT/_0217_ ), .B2(\CLINT/_0365_ ), .ZN(\CLINT/_0040_ ) );
AND2_X1 \CLINT/_1045_ ( .A1(\CLINT/_0217_ ), .A2(\CLINT/_0228_ ), .ZN(\CLINT/_0368_ ) );
AND2_X1 \CLINT/_1046_ ( .A1(\CLINT/_0365_ ), .A2(\CLINT/_0368_ ), .ZN(\CLINT/_0369_ ) );
AOI21_X1 \CLINT/_1047_ ( .A(\CLINT/_0228_ ), .B1(\CLINT/_0365_ ), .B2(\CLINT/_0217_ ), .ZN(\CLINT/_0370_ ) );
NOR3_X1 \CLINT/_1048_ ( .A1(\CLINT/_0369_ ), .A2(\CLINT/_0370_ ), .A3(fanout_net_7 ), .ZN(\CLINT/_0041_ ) );
OAI21_X1 \CLINT/_1049_ ( .A(\CLINT/_0358_ ), .B1(\CLINT/_0369_ ), .B2(\CLINT/_0233_ ), .ZN(\CLINT/_0371_ ) );
AOI21_X1 \CLINT/_1050_ ( .A(\CLINT/_0371_ ), .B1(\CLINT/_0233_ ), .B2(\CLINT/_0369_ ), .ZN(\CLINT/_0042_ ) );
AOI21_X1 \CLINT/_1051_ ( .A(\CLINT/_0234_ ), .B1(\CLINT/_0369_ ), .B2(\CLINT/_0233_ ), .ZN(\CLINT/_0372_ ) );
AND4_X1 \CLINT/_1052_ ( .A1(\CLINT/_0217_ ), .A2(\CLINT/_0228_ ), .A3(\CLINT/_0233_ ), .A4(\CLINT/_0234_ ), .ZN(\CLINT/_0373_ ) );
AND2_X4 \CLINT/_1053_ ( .A1(\CLINT/_0365_ ), .A2(\CLINT/_0373_ ), .ZN(\CLINT/_0374_ ) );
NOR3_X1 \CLINT/_1054_ ( .A1(\CLINT/_0372_ ), .A2(fanout_net_7 ), .A3(\CLINT/_0374_ ), .ZN(\CLINT/_0043_ ) );
AND4_X2 \CLINT/_1055_ ( .A1(\CLINT/_0195_ ), .A2(\CLINT/_0206_ ), .A3(\CLINT/_0228_ ), .A4(\CLINT/_0233_ ), .ZN(\CLINT/_0375_ ) );
AND4_X2 \CLINT/_1056_ ( .A1(\CLINT/_0173_ ), .A2(\CLINT/_0184_ ), .A3(\CLINT/_0217_ ), .A4(\CLINT/_0234_ ), .ZN(\CLINT/_0376_ ) );
AND2_X4 \CLINT/_1057_ ( .A1(\CLINT/_0375_ ), .A2(\CLINT/_0376_ ), .ZN(\CLINT/_0377_ ) );
OAI21_X1 \CLINT/_1058_ ( .A(\CLINT/_0358_ ), .B1(\CLINT/_0377_ ), .B2(\CLINT/_0235_ ), .ZN(\CLINT/_0378_ ) );
AOI21_X1 \CLINT/_1059_ ( .A(\CLINT/_0378_ ), .B1(\CLINT/_0235_ ), .B2(\CLINT/_0377_ ), .ZN(\CLINT/_0044_ ) );
AOI21_X1 \CLINT/_1060_ ( .A(\CLINT/_0236_ ), .B1(\CLINT/_0377_ ), .B2(\CLINT/_0235_ ), .ZN(\CLINT/_0379_ ) );
AND2_X4 \CLINT/_1061_ ( .A1(\CLINT/_0235_ ), .A2(\CLINT/_0236_ ), .ZN(\CLINT/_0380_ ) );
AOI211_X4 \CLINT/_1062_ ( .A(fanout_net_7 ), .B(\CLINT/_0379_ ), .C1(\CLINT/_0374_ ), .C2(\CLINT/_0380_ ), .ZN(\CLINT/_0045_ ) );
AND2_X1 \CLINT/_1063_ ( .A1(\CLINT/_0374_ ), .A2(\CLINT/_0380_ ), .ZN(\CLINT/_0381_ ) );
OAI21_X1 \CLINT/_1064_ ( .A(\CLINT/_0358_ ), .B1(\CLINT/_0381_ ), .B2(\CLINT/_0174_ ), .ZN(\CLINT/_0382_ ) );
AOI21_X1 \CLINT/_1065_ ( .A(\CLINT/_0382_ ), .B1(\CLINT/_0174_ ), .B2(\CLINT/_0381_ ), .ZN(\CLINT/_0046_ ) );
AND2_X4 \CLINT/_1066_ ( .A1(\CLINT/_0174_ ), .A2(\CLINT/_0175_ ), .ZN(\CLINT/_0383_ ) );
AND2_X1 \CLINT/_1067_ ( .A1(\CLINT/_0381_ ), .A2(\CLINT/_0383_ ), .ZN(\CLINT/_0384_ ) );
AOI21_X1 \CLINT/_1068_ ( .A(\CLINT/_0175_ ), .B1(\CLINT/_0381_ ), .B2(\CLINT/_0174_ ), .ZN(\CLINT/_0385_ ) );
NOR3_X1 \CLINT/_1069_ ( .A1(\CLINT/_0384_ ), .A2(\CLINT/_0385_ ), .A3(fanout_net_7 ), .ZN(\CLINT/_0047_ ) );
AND2_X4 \CLINT/_1070_ ( .A1(\CLINT/_0380_ ), .A2(\CLINT/_0383_ ), .ZN(\CLINT/_0386_ ) );
AND3_X1 \CLINT/_1071_ ( .A1(\CLINT/_0386_ ), .A2(\CLINT/_0375_ ), .A3(\CLINT/_0376_ ), .ZN(\CLINT/_0387_ ) );
OAI21_X1 \CLINT/_1072_ ( .A(\CLINT/_0359_ ), .B1(\CLINT/_0387_ ), .B2(\CLINT/_0176_ ), .ZN(\CLINT/_0388_ ) );
AND3_X1 \CLINT/_1073_ ( .A1(\CLINT/_0377_ ), .A2(\CLINT/_0176_ ), .A3(\CLINT/_0386_ ), .ZN(\CLINT/_0389_ ) );
NOR2_X1 \CLINT/_1074_ ( .A1(\CLINT/_0388_ ), .A2(\CLINT/_0389_ ), .ZN(\CLINT/_0048_ ) );
AND3_X1 \CLINT/_1075_ ( .A1(\CLINT/_0387_ ), .A2(\CLINT/_0176_ ), .A3(\CLINT/_0177_ ), .ZN(\CLINT/_0390_ ) );
AOI21_X1 \CLINT/_1076_ ( .A(\CLINT/_0177_ ), .B1(\CLINT/_0387_ ), .B2(\CLINT/_0176_ ), .ZN(\CLINT/_0391_ ) );
NOR3_X1 \CLINT/_1077_ ( .A1(\CLINT/_0390_ ), .A2(\CLINT/_0391_ ), .A3(fanout_net_7 ), .ZN(\CLINT/_0049_ ) );
OAI21_X1 \CLINT/_1078_ ( .A(\CLINT/_0359_ ), .B1(\CLINT/_0390_ ), .B2(\CLINT/_0178_ ), .ZN(\CLINT/_0392_ ) );
AND3_X1 \CLINT/_1079_ ( .A1(\CLINT/_0389_ ), .A2(\CLINT/_0177_ ), .A3(\CLINT/_0178_ ), .ZN(\CLINT/_0393_ ) );
NOR2_X1 \CLINT/_1080_ ( .A1(\CLINT/_0392_ ), .A2(\CLINT/_0393_ ), .ZN(\CLINT/_0050_ ) );
AOI21_X1 \CLINT/_1081_ ( .A(\CLINT/_0179_ ), .B1(\CLINT/_0390_ ), .B2(\CLINT/_0178_ ), .ZN(\CLINT/_0394_ ) );
AND4_X1 \CLINT/_1082_ ( .A1(\CLINT/_0177_ ), .A2(\CLINT/_0389_ ), .A3(\CLINT/_0178_ ), .A4(\CLINT/_0179_ ), .ZN(\CLINT/_0395_ ) );
NOR3_X1 \CLINT/_1083_ ( .A1(\CLINT/_0394_ ), .A2(\CLINT/_0395_ ), .A3(fanout_net_7 ), .ZN(\CLINT/_0051_ ) );
AND2_X4 \CLINT/_1084_ ( .A1(\CLINT/_0178_ ), .A2(\CLINT/_0179_ ), .ZN(\CLINT/_0396_ ) );
AND3_X2 \CLINT/_1085_ ( .A1(\CLINT/_0396_ ), .A2(\CLINT/_0176_ ), .A3(\CLINT/_0177_ ), .ZN(\CLINT/_0397_ ) );
AND2_X4 \CLINT/_1086_ ( .A1(\CLINT/_0397_ ), .A2(\CLINT/_0386_ ), .ZN(\CLINT/_0398_ ) );
AND2_X4 \CLINT/_1087_ ( .A1(\CLINT/_0398_ ), .A2(\CLINT/_0377_ ), .ZN(\CLINT/_0399_ ) );
OAI21_X1 \CLINT/_1088_ ( .A(\CLINT/_0359_ ), .B1(\CLINT/_0399_ ), .B2(\CLINT/_0180_ ), .ZN(\CLINT/_0400_ ) );
AND3_X1 \CLINT/_1089_ ( .A1(\CLINT/_0398_ ), .A2(\CLINT/_0180_ ), .A3(\CLINT/_0377_ ), .ZN(\CLINT/_0401_ ) );
NOR2_X1 \CLINT/_1090_ ( .A1(\CLINT/_0400_ ), .A2(\CLINT/_0401_ ), .ZN(\CLINT/_0052_ ) );
AND2_X1 \CLINT/_1091_ ( .A1(\CLINT/_0401_ ), .A2(\CLINT/_0181_ ), .ZN(\CLINT/_0402_ ) );
NOR2_X1 \CLINT/_1092_ ( .A1(\CLINT/_0401_ ), .A2(\CLINT/_0181_ ), .ZN(\CLINT/_0403_ ) );
NOR3_X1 \CLINT/_1093_ ( .A1(\CLINT/_0402_ ), .A2(\CLINT/_0403_ ), .A3(fanout_net_7 ), .ZN(\CLINT/_0053_ ) );
OAI21_X1 \CLINT/_1094_ ( .A(\CLINT/_0359_ ), .B1(\CLINT/_0402_ ), .B2(\CLINT/_0182_ ), .ZN(\CLINT/_0404_ ) );
AND3_X1 \CLINT/_1095_ ( .A1(\CLINT/_0401_ ), .A2(\CLINT/_0181_ ), .A3(\CLINT/_0182_ ), .ZN(\CLINT/_0405_ ) );
NOR2_X1 \CLINT/_1096_ ( .A1(\CLINT/_0404_ ), .A2(\CLINT/_0405_ ), .ZN(\CLINT/_0054_ ) );
NOR2_X1 \CLINT/_1097_ ( .A1(\CLINT/_0405_ ), .A2(\CLINT/_0183_ ), .ZN(\CLINT/_0406_ ) );
AND2_X1 \CLINT/_1098_ ( .A1(\CLINT/_0374_ ), .A2(\CLINT/_0398_ ), .ZN(\CLINT/_0407_ ) );
AND2_X4 \CLINT/_1099_ ( .A1(\CLINT/_0180_ ), .A2(\CLINT/_0181_ ), .ZN(\CLINT/_0408_ ) );
AND2_X4 \CLINT/_1100_ ( .A1(\CLINT/_0182_ ), .A2(\CLINT/_0183_ ), .ZN(\CLINT/_0409_ ) );
AND2_X4 \CLINT/_1101_ ( .A1(\CLINT/_0408_ ), .A2(\CLINT/_0409_ ), .ZN(\CLINT/_0410_ ) );
AND2_X1 \CLINT/_1102_ ( .A1(\CLINT/_0407_ ), .A2(\CLINT/_0410_ ), .ZN(\CLINT/_0411_ ) );
NOR3_X1 \CLINT/_1103_ ( .A1(\CLINT/_0406_ ), .A2(\CLINT/_0411_ ), .A3(fanout_net_7 ), .ZN(\CLINT/_0055_ ) );
AND3_X1 \CLINT/_1104_ ( .A1(\CLINT/_0398_ ), .A2(\CLINT/_0377_ ), .A3(\CLINT/_0410_ ), .ZN(\CLINT/_0412_ ) );
AND2_X1 \CLINT/_1105_ ( .A1(\CLINT/_0412_ ), .A2(\CLINT/_0185_ ), .ZN(\CLINT/_0413_ ) );
OAI21_X1 \CLINT/_1106_ ( .A(\CLINT/_0363_ ), .B1(\CLINT/_0412_ ), .B2(\CLINT/_0185_ ), .ZN(\CLINT/_0414_ ) );
NOR2_X1 \CLINT/_1107_ ( .A1(\CLINT/_0413_ ), .A2(\CLINT/_0414_ ), .ZN(\CLINT/_0056_ ) );
AND3_X1 \CLINT/_1108_ ( .A1(\CLINT/_0412_ ), .A2(\CLINT/_0185_ ), .A3(\CLINT/_0186_ ), .ZN(\CLINT/_0415_ ) );
AOI21_X1 \CLINT/_1109_ ( .A(\CLINT/_0186_ ), .B1(\CLINT/_0412_ ), .B2(\CLINT/_0185_ ), .ZN(\CLINT/_0416_ ) );
NOR3_X1 \CLINT/_1110_ ( .A1(\CLINT/_0415_ ), .A2(\CLINT/_0416_ ), .A3(fanout_net_7 ), .ZN(\CLINT/_0057_ ) );
AND2_X1 \CLINT/_1111_ ( .A1(\CLINT/_0415_ ), .A2(\CLINT/_0187_ ), .ZN(\CLINT/_0417_ ) );
OAI21_X1 \CLINT/_1112_ ( .A(\CLINT/_0363_ ), .B1(\CLINT/_0415_ ), .B2(\CLINT/_0187_ ), .ZN(\CLINT/_0418_ ) );
NOR2_X1 \CLINT/_1113_ ( .A1(\CLINT/_0417_ ), .A2(\CLINT/_0418_ ), .ZN(\CLINT/_0058_ ) );
AND3_X1 \CLINT/_1114_ ( .A1(\CLINT/_0415_ ), .A2(\CLINT/_0187_ ), .A3(\CLINT/_0188_ ), .ZN(\CLINT/_0419_ ) );
AOI21_X1 \CLINT/_1115_ ( .A(\CLINT/_0188_ ), .B1(\CLINT/_0415_ ), .B2(\CLINT/_0187_ ), .ZN(\CLINT/_0420_ ) );
NOR3_X1 \CLINT/_1116_ ( .A1(\CLINT/_0419_ ), .A2(\CLINT/_0420_ ), .A3(fanout_net_7 ), .ZN(\CLINT/_0059_ ) );
AND2_X4 \CLINT/_1117_ ( .A1(\CLINT/_0185_ ), .A2(\CLINT/_0186_ ), .ZN(\CLINT/_0421_ ) );
AND2_X4 \CLINT/_1118_ ( .A1(\CLINT/_0187_ ), .A2(\CLINT/_0188_ ), .ZN(\CLINT/_0422_ ) );
AND2_X1 \CLINT/_1119_ ( .A1(\CLINT/_0421_ ), .A2(\CLINT/_0422_ ), .ZN(\CLINT/_0423_ ) );
AND2_X1 \CLINT/_1120_ ( .A1(\CLINT/_0412_ ), .A2(\CLINT/_0423_ ), .ZN(\CLINT/_0424_ ) );
OAI21_X1 \CLINT/_1121_ ( .A(\CLINT/_0359_ ), .B1(\CLINT/_0424_ ), .B2(\CLINT/_0189_ ), .ZN(\CLINT/_0425_ ) );
AND3_X1 \CLINT/_1122_ ( .A1(\CLINT/_0412_ ), .A2(\CLINT/_0189_ ), .A3(\CLINT/_0423_ ), .ZN(\CLINT/_0426_ ) );
NOR2_X1 \CLINT/_1123_ ( .A1(\CLINT/_0425_ ), .A2(\CLINT/_0426_ ), .ZN(\CLINT/_0060_ ) );
AND2_X1 \CLINT/_1124_ ( .A1(\CLINT/_0426_ ), .A2(\CLINT/_0190_ ), .ZN(\CLINT/_0427_ ) );
NOR2_X1 \CLINT/_1125_ ( .A1(\CLINT/_0426_ ), .A2(\CLINT/_0190_ ), .ZN(\CLINT/_0428_ ) );
NOR3_X1 \CLINT/_1126_ ( .A1(\CLINT/_0427_ ), .A2(\CLINT/_0428_ ), .A3(fanout_net_7 ), .ZN(\CLINT/_0061_ ) );
OAI21_X1 \CLINT/_1127_ ( .A(\CLINT/_0359_ ), .B1(\CLINT/_0427_ ), .B2(\CLINT/_0191_ ), .ZN(\CLINT/_0429_ ) );
AND3_X1 \CLINT/_1128_ ( .A1(\CLINT/_0426_ ), .A2(\CLINT/_0190_ ), .A3(\CLINT/_0191_ ), .ZN(\CLINT/_0430_ ) );
NOR2_X1 \CLINT/_1129_ ( .A1(\CLINT/_0429_ ), .A2(\CLINT/_0430_ ), .ZN(\CLINT/_0062_ ) );
AOI21_X1 \CLINT/_1130_ ( .A(\CLINT/_0192_ ), .B1(\CLINT/_0427_ ), .B2(\CLINT/_0191_ ), .ZN(\CLINT/_0431_ ) );
AND4_X1 \CLINT/_1131_ ( .A1(\CLINT/_0190_ ), .A2(\CLINT/_0426_ ), .A3(\CLINT/_0191_ ), .A4(\CLINT/_0192_ ), .ZN(\CLINT/_0432_ ) );
NOR3_X1 \CLINT/_1132_ ( .A1(\CLINT/_0431_ ), .A2(\CLINT/_0432_ ), .A3(fanout_net_7 ), .ZN(\CLINT/_0063_ ) );
NAND2_X4 \CLINT/_1133_ ( .A1(\CLINT/_0190_ ), .A2(\CLINT/_0191_ ), .ZN(\CLINT/_0433_ ) );
NAND2_X4 \CLINT/_1134_ ( .A1(\CLINT/_0189_ ), .A2(\CLINT/_0192_ ), .ZN(\CLINT/_0434_ ) );
NOR2_X4 \CLINT/_1135_ ( .A1(\CLINT/_0433_ ), .A2(\CLINT/_0434_ ), .ZN(\CLINT/_0435_ ) );
AND3_X1 \CLINT/_1136_ ( .A1(\CLINT/_0412_ ), .A2(\CLINT/_0423_ ), .A3(\CLINT/_0435_ ), .ZN(\CLINT/_0436_ ) );
AND2_X1 \CLINT/_1137_ ( .A1(\CLINT/_0436_ ), .A2(\CLINT/_0193_ ), .ZN(\CLINT/_0437_ ) );
OAI21_X1 \CLINT/_1138_ ( .A(\CLINT/_0363_ ), .B1(\CLINT/_0436_ ), .B2(\CLINT/_0193_ ), .ZN(\CLINT/_0438_ ) );
NOR2_X1 \CLINT/_1139_ ( .A1(\CLINT/_0437_ ), .A2(\CLINT/_0438_ ), .ZN(\CLINT/_0064_ ) );
AND3_X1 \CLINT/_1140_ ( .A1(\CLINT/_0436_ ), .A2(\CLINT/_0193_ ), .A3(\CLINT/_0194_ ), .ZN(\CLINT/_0439_ ) );
AOI21_X1 \CLINT/_1141_ ( .A(\CLINT/_0194_ ), .B1(\CLINT/_0436_ ), .B2(\CLINT/_0193_ ), .ZN(\CLINT/_0440_ ) );
NOR3_X1 \CLINT/_1142_ ( .A1(\CLINT/_0439_ ), .A2(\CLINT/_0440_ ), .A3(fanout_net_7 ), .ZN(\CLINT/_0065_ ) );
AND2_X1 \CLINT/_1143_ ( .A1(\CLINT/_0439_ ), .A2(\CLINT/_0196_ ), .ZN(\CLINT/_0441_ ) );
OAI21_X1 \CLINT/_1144_ ( .A(\CLINT/_0363_ ), .B1(\CLINT/_0439_ ), .B2(\CLINT/_0196_ ), .ZN(\CLINT/_0442_ ) );
NOR2_X1 \CLINT/_1145_ ( .A1(\CLINT/_0441_ ), .A2(\CLINT/_0442_ ), .ZN(\CLINT/_0066_ ) );
AOI21_X1 \CLINT/_1146_ ( .A(\CLINT/_0197_ ), .B1(\CLINT/_0439_ ), .B2(\CLINT/_0196_ ), .ZN(\CLINT/_0443_ ) );
INV_X1 \CLINT/_1147_ ( .A(\CLINT/_0407_ ), .ZN(\CLINT/_0444_ ) );
INV_X4 \CLINT/_1148_ ( .A(\CLINT/_0410_ ), .ZN(\CLINT/_0445_ ) );
AND3_X4 \CLINT/_1149_ ( .A1(\CLINT/_0435_ ), .A2(\CLINT/_0421_ ), .A3(\CLINT/_0422_ ), .ZN(\CLINT/_0446_ ) );
INV_X2 \CLINT/_1150_ ( .A(\CLINT/_0446_ ), .ZN(\CLINT/_0447_ ) );
AND2_X1 \CLINT/_1151_ ( .A1(\CLINT/_0193_ ), .A2(\CLINT/_0197_ ), .ZN(\CLINT/_0448_ ) );
NAND3_X4 \CLINT/_1152_ ( .A1(\CLINT/_0448_ ), .A2(\CLINT/_0194_ ), .A3(\CLINT/_0196_ ), .ZN(\CLINT/_0449_ ) );
NOR4_X1 \CLINT/_1153_ ( .A1(\CLINT/_0444_ ), .A2(\CLINT/_0445_ ), .A3(\CLINT/_0447_ ), .A4(\CLINT/_0449_ ), .ZN(\CLINT/_0450_ ) );
NOR3_X1 \CLINT/_1154_ ( .A1(\CLINT/_0443_ ), .A2(fanout_net_7 ), .A3(\CLINT/_0450_ ), .ZN(\CLINT/_0067_ ) );
NOR3_X4 \CLINT/_1155_ ( .A1(\CLINT/_0447_ ), .A2(\CLINT/_0449_ ), .A3(\CLINT/_0445_ ), .ZN(\CLINT/_0451_ ) );
AND2_X4 \CLINT/_1156_ ( .A1(\CLINT/_0451_ ), .A2(\CLINT/_0399_ ), .ZN(\CLINT/_0452_ ) );
OAI21_X1 \CLINT/_1157_ ( .A(\CLINT/_0359_ ), .B1(\CLINT/_0452_ ), .B2(\CLINT/_0198_ ), .ZN(\CLINT/_0453_ ) );
AND3_X1 \CLINT/_1158_ ( .A1(\CLINT/_0451_ ), .A2(\CLINT/_0198_ ), .A3(\CLINT/_0399_ ), .ZN(\CLINT/_0454_ ) );
NOR2_X1 \CLINT/_1159_ ( .A1(\CLINT/_0453_ ), .A2(\CLINT/_0454_ ), .ZN(\CLINT/_0068_ ) );
NAND3_X1 \CLINT/_1160_ ( .A1(\CLINT/_0451_ ), .A2(\CLINT/_0399_ ), .A3(\CLINT/_0198_ ), .ZN(\CLINT/_0455_ ) );
XNOR2_X1 \CLINT/_1161_ ( .A(\CLINT/_0455_ ), .B(\CLINT/_0199_ ), .ZN(\CLINT/_0456_ ) );
AND2_X1 \CLINT/_1162_ ( .A1(\CLINT/_0456_ ), .A2(\CLINT/_0359_ ), .ZN(\CLINT/_0069_ ) );
AND2_X4 \CLINT/_1163_ ( .A1(\CLINT/_0198_ ), .A2(\CLINT/_0199_ ), .ZN(\CLINT/_0457_ ) );
AND3_X1 \CLINT/_1164_ ( .A1(\CLINT/_0407_ ), .A2(\CLINT/_0451_ ), .A3(\CLINT/_0457_ ), .ZN(\CLINT/_0458_ ) );
OAI21_X1 \CLINT/_1165_ ( .A(\CLINT/_0363_ ), .B1(\CLINT/_0458_ ), .B2(\CLINT/_0200_ ), .ZN(\CLINT/_0459_ ) );
AND3_X1 \CLINT/_1166_ ( .A1(\CLINT/_0454_ ), .A2(\CLINT/_0199_ ), .A3(\CLINT/_0200_ ), .ZN(\CLINT/_0460_ ) );
NOR2_X1 \CLINT/_1167_ ( .A1(\CLINT/_0459_ ), .A2(\CLINT/_0460_ ), .ZN(\CLINT/_0070_ ) );
AOI21_X1 \CLINT/_1168_ ( .A(\CLINT/_0201_ ), .B1(\CLINT/_0458_ ), .B2(\CLINT/_0200_ ), .ZN(\CLINT/_0461_ ) );
AND4_X1 \CLINT/_1169_ ( .A1(\CLINT/_0199_ ), .A2(\CLINT/_0454_ ), .A3(\CLINT/_0200_ ), .A4(\CLINT/_0201_ ), .ZN(\CLINT/_0462_ ) );
NOR3_X1 \CLINT/_1170_ ( .A1(\CLINT/_0461_ ), .A2(\CLINT/_0462_ ), .A3(fanout_net_7 ), .ZN(\CLINT/_0071_ ) );
AND2_X4 \CLINT/_1171_ ( .A1(\CLINT/_0200_ ), .A2(\CLINT/_0201_ ), .ZN(\CLINT/_0463_ ) );
AND2_X4 \CLINT/_1172_ ( .A1(\CLINT/_0457_ ), .A2(\CLINT/_0463_ ), .ZN(\CLINT/_0464_ ) );
AND3_X1 \CLINT/_1173_ ( .A1(\CLINT/_0451_ ), .A2(\CLINT/_0399_ ), .A3(\CLINT/_0464_ ), .ZN(\CLINT/_0465_ ) );
AND2_X1 \CLINT/_1174_ ( .A1(\CLINT/_0465_ ), .A2(\CLINT/_0202_ ), .ZN(\CLINT/_0466_ ) );
BUF_X4 \CLINT/_1175_ ( .A(\CLINT/_0358_ ), .Z(\CLINT/_0467_ ) );
OAI21_X1 \CLINT/_1176_ ( .A(\CLINT/_0467_ ), .B1(\CLINT/_0465_ ), .B2(\CLINT/_0202_ ), .ZN(\CLINT/_0468_ ) );
NOR2_X1 \CLINT/_1177_ ( .A1(\CLINT/_0466_ ), .A2(\CLINT/_0468_ ), .ZN(\CLINT/_0072_ ) );
AND3_X1 \CLINT/_1178_ ( .A1(\CLINT/_0465_ ), .A2(\CLINT/_0202_ ), .A3(\CLINT/_0203_ ), .ZN(\CLINT/_0469_ ) );
AOI21_X1 \CLINT/_1179_ ( .A(\CLINT/_0203_ ), .B1(\CLINT/_0465_ ), .B2(\CLINT/_0202_ ), .ZN(\CLINT/_0470_ ) );
NOR3_X1 \CLINT/_1180_ ( .A1(\CLINT/_0469_ ), .A2(\CLINT/_0470_ ), .A3(fanout_net_7 ), .ZN(\CLINT/_0073_ ) );
AND2_X1 \CLINT/_1181_ ( .A1(\CLINT/_0469_ ), .A2(\CLINT/_0204_ ), .ZN(\CLINT/_0471_ ) );
OAI21_X1 \CLINT/_1182_ ( .A(\CLINT/_0467_ ), .B1(\CLINT/_0469_ ), .B2(\CLINT/_0204_ ), .ZN(\CLINT/_0472_ ) );
NOR2_X1 \CLINT/_1183_ ( .A1(\CLINT/_0471_ ), .A2(\CLINT/_0472_ ), .ZN(\CLINT/_0074_ ) );
AOI21_X1 \CLINT/_1184_ ( .A(\CLINT/_0205_ ), .B1(\CLINT/_0469_ ), .B2(\CLINT/_0204_ ), .ZN(\CLINT/_0473_ ) );
AND2_X1 \CLINT/_1185_ ( .A1(\CLINT/_0407_ ), .A2(\CLINT/_0451_ ), .ZN(\CLINT/_0474_ ) );
AND4_X4 \CLINT/_1186_ ( .A1(\CLINT/_0202_ ), .A2(\CLINT/_0203_ ), .A3(\CLINT/_0204_ ), .A4(\CLINT/_0205_ ), .ZN(\CLINT/_0475_ ) );
AND2_X1 \CLINT/_1187_ ( .A1(\CLINT/_0464_ ), .A2(\CLINT/_0475_ ), .ZN(\CLINT/_0476_ ) );
AND2_X1 \CLINT/_1188_ ( .A1(\CLINT/_0474_ ), .A2(\CLINT/_0476_ ), .ZN(\CLINT/_0477_ ) );
NOR3_X1 \CLINT/_1189_ ( .A1(\CLINT/_0473_ ), .A2(fanout_net_7 ), .A3(\CLINT/_0477_ ), .ZN(\CLINT/_0075_ ) );
AND3_X1 \CLINT/_1190_ ( .A1(\CLINT/_0451_ ), .A2(\CLINT/_0399_ ), .A3(\CLINT/_0476_ ), .ZN(\CLINT/_0478_ ) );
AND2_X1 \CLINT/_1191_ ( .A1(\CLINT/_0478_ ), .A2(\CLINT/_0207_ ), .ZN(\CLINT/_0479_ ) );
OAI21_X1 \CLINT/_1192_ ( .A(\CLINT/_0467_ ), .B1(\CLINT/_0478_ ), .B2(\CLINT/_0207_ ), .ZN(\CLINT/_0480_ ) );
NOR2_X1 \CLINT/_1193_ ( .A1(\CLINT/_0479_ ), .A2(\CLINT/_0480_ ), .ZN(\CLINT/_0076_ ) );
AND3_X1 \CLINT/_1194_ ( .A1(\CLINT/_0478_ ), .A2(\CLINT/_0207_ ), .A3(\CLINT/_0208_ ), .ZN(\CLINT/_0481_ ) );
AOI21_X1 \CLINT/_1195_ ( .A(\CLINT/_0208_ ), .B1(\CLINT/_0478_ ), .B2(\CLINT/_0207_ ), .ZN(\CLINT/_0482_ ) );
NOR3_X1 \CLINT/_1196_ ( .A1(\CLINT/_0481_ ), .A2(\CLINT/_0482_ ), .A3(fanout_net_7 ), .ZN(\CLINT/_0077_ ) );
AND2_X1 \CLINT/_1197_ ( .A1(\CLINT/_0481_ ), .A2(\CLINT/_0209_ ), .ZN(\CLINT/_0483_ ) );
OAI21_X1 \CLINT/_1198_ ( .A(\CLINT/_0467_ ), .B1(\CLINT/_0481_ ), .B2(\CLINT/_0209_ ), .ZN(\CLINT/_0484_ ) );
NOR2_X1 \CLINT/_1199_ ( .A1(\CLINT/_0483_ ), .A2(\CLINT/_0484_ ), .ZN(\CLINT/_0078_ ) );
AOI21_X1 \CLINT/_1200_ ( .A(\CLINT/_0210_ ), .B1(\CLINT/_0481_ ), .B2(\CLINT/_0209_ ), .ZN(\CLINT/_0485_ ) );
NAND2_X1 \CLINT/_1201_ ( .A1(\CLINT/_0208_ ), .A2(\CLINT/_0209_ ), .ZN(\CLINT/_0486_ ) );
NAND2_X1 \CLINT/_1202_ ( .A1(\CLINT/_0207_ ), .A2(\CLINT/_0210_ ), .ZN(\CLINT/_0487_ ) );
NOR2_X1 \CLINT/_1203_ ( .A1(\CLINT/_0486_ ), .A2(\CLINT/_0487_ ), .ZN(\CLINT/_0488_ ) );
AND2_X1 \CLINT/_1204_ ( .A1(\CLINT/_0478_ ), .A2(\CLINT/_0488_ ), .ZN(\CLINT/_0489_ ) );
NOR3_X1 \CLINT/_1205_ ( .A1(\CLINT/_0485_ ), .A2(fanout_net_7 ), .A3(\CLINT/_0489_ ), .ZN(\CLINT/_0079_ ) );
OAI21_X1 \CLINT/_1206_ ( .A(\CLINT/_0363_ ), .B1(\CLINT/_0489_ ), .B2(\CLINT/_0211_ ), .ZN(\CLINT/_0490_ ) );
AND3_X1 \CLINT/_1207_ ( .A1(\CLINT/_0478_ ), .A2(\CLINT/_0211_ ), .A3(\CLINT/_0488_ ), .ZN(\CLINT/_0491_ ) );
NOR2_X1 \CLINT/_1208_ ( .A1(\CLINT/_0490_ ), .A2(\CLINT/_0491_ ), .ZN(\CLINT/_0080_ ) );
AND2_X1 \CLINT/_1209_ ( .A1(\CLINT/_0491_ ), .A2(\CLINT/_0212_ ), .ZN(\CLINT/_0492_ ) );
NOR2_X1 \CLINT/_1210_ ( .A1(\CLINT/_0491_ ), .A2(\CLINT/_0212_ ), .ZN(\CLINT/_0493_ ) );
NOR3_X1 \CLINT/_1211_ ( .A1(\CLINT/_0492_ ), .A2(\CLINT/_0493_ ), .A3(fanout_net_7 ), .ZN(\CLINT/_0081_ ) );
OAI21_X1 \CLINT/_1212_ ( .A(\CLINT/_0363_ ), .B1(\CLINT/_0492_ ), .B2(\CLINT/_0213_ ), .ZN(\CLINT/_0494_ ) );
AND3_X2 \CLINT/_1213_ ( .A1(\CLINT/_0491_ ), .A2(\CLINT/_0212_ ), .A3(\CLINT/_0213_ ), .ZN(\CLINT/_0495_ ) );
NOR2_X1 \CLINT/_1214_ ( .A1(\CLINT/_0494_ ), .A2(\CLINT/_0495_ ), .ZN(\CLINT/_0082_ ) );
NOR2_X1 \CLINT/_1215_ ( .A1(\CLINT/_0495_ ), .A2(\CLINT/_0214_ ), .ZN(\CLINT/_0496_ ) );
AND2_X1 \CLINT/_1216_ ( .A1(\CLINT/_0211_ ), .A2(\CLINT/_0214_ ), .ZN(\CLINT/_0497_ ) );
AND3_X1 \CLINT/_1217_ ( .A1(\CLINT/_0497_ ), .A2(\CLINT/_0212_ ), .A3(\CLINT/_0213_ ), .ZN(\CLINT/_0498_ ) );
AND4_X1 \CLINT/_1218_ ( .A1(\CLINT/_0474_ ), .A2(\CLINT/_0476_ ), .A3(\CLINT/_0488_ ), .A4(\CLINT/_0498_ ), .ZN(\CLINT/_0499_ ) );
NOR3_X1 \CLINT/_1219_ ( .A1(\CLINT/_0496_ ), .A2(fanout_net_7 ), .A3(\CLINT/_0499_ ), .ZN(\CLINT/_0083_ ) );
AND3_X1 \CLINT/_1220_ ( .A1(\CLINT/_0476_ ), .A2(\CLINT/_0488_ ), .A3(\CLINT/_0498_ ), .ZN(\CLINT/_0500_ ) );
AND2_X1 \CLINT/_1221_ ( .A1(\CLINT/_0452_ ), .A2(\CLINT/_0500_ ), .ZN(\CLINT/_0501_ ) );
OAI21_X1 \CLINT/_1222_ ( .A(\CLINT/_0363_ ), .B1(\CLINT/_0501_ ), .B2(\CLINT/_0215_ ), .ZN(\CLINT/_0502_ ) );
AND3_X1 \CLINT/_1223_ ( .A1(\CLINT/_0452_ ), .A2(\CLINT/_0215_ ), .A3(\CLINT/_0500_ ), .ZN(\CLINT/_0503_ ) );
NOR2_X1 \CLINT/_1224_ ( .A1(\CLINT/_0502_ ), .A2(\CLINT/_0503_ ), .ZN(\CLINT/_0084_ ) );
NAND3_X1 \CLINT/_1225_ ( .A1(\CLINT/_0452_ ), .A2(\CLINT/_0215_ ), .A3(\CLINT/_0500_ ), .ZN(\CLINT/_0504_ ) );
XNOR2_X1 \CLINT/_1226_ ( .A(\CLINT/_0504_ ), .B(\CLINT/_0216_ ), .ZN(\CLINT/_0505_ ) );
AND2_X1 \CLINT/_1227_ ( .A1(\CLINT/_0505_ ), .A2(\CLINT/_0359_ ), .ZN(\CLINT/_0085_ ) );
AND2_X1 \CLINT/_1228_ ( .A1(\CLINT/_0215_ ), .A2(\CLINT/_0216_ ), .ZN(\CLINT/_0506_ ) );
AND3_X1 \CLINT/_1229_ ( .A1(\CLINT/_0474_ ), .A2(\CLINT/_0500_ ), .A3(\CLINT/_0506_ ), .ZN(\CLINT/_0507_ ) );
OAI21_X1 \CLINT/_1230_ ( .A(\CLINT/_0363_ ), .B1(\CLINT/_0507_ ), .B2(\CLINT/_0218_ ), .ZN(\CLINT/_0508_ ) );
AND3_X1 \CLINT/_1231_ ( .A1(\CLINT/_0503_ ), .A2(\CLINT/_0216_ ), .A3(\CLINT/_0218_ ), .ZN(\CLINT/_0509_ ) );
NOR2_X1 \CLINT/_1232_ ( .A1(\CLINT/_0508_ ), .A2(\CLINT/_0509_ ), .ZN(\CLINT/_0086_ ) );
AOI21_X1 \CLINT/_1233_ ( .A(\CLINT/_0219_ ), .B1(\CLINT/_0507_ ), .B2(\CLINT/_0218_ ), .ZN(\CLINT/_0510_ ) );
AND4_X1 \CLINT/_1234_ ( .A1(\CLINT/_0216_ ), .A2(\CLINT/_0503_ ), .A3(\CLINT/_0218_ ), .A4(\CLINT/_0219_ ), .ZN(\CLINT/_0511_ ) );
NOR3_X1 \CLINT/_1235_ ( .A1(\CLINT/_0510_ ), .A2(\CLINT/_0511_ ), .A3(fanout_net_7 ), .ZN(\CLINT/_0087_ ) );
AND2_X1 \CLINT/_1236_ ( .A1(\CLINT/_0218_ ), .A2(\CLINT/_0219_ ), .ZN(\CLINT/_0512_ ) );
AND2_X1 \CLINT/_1237_ ( .A1(\CLINT/_0506_ ), .A2(\CLINT/_0512_ ), .ZN(\CLINT/_0513_ ) );
AND3_X1 \CLINT/_1238_ ( .A1(\CLINT/_0452_ ), .A2(\CLINT/_0500_ ), .A3(\CLINT/_0513_ ), .ZN(\CLINT/_0514_ ) );
AND2_X1 \CLINT/_1239_ ( .A1(\CLINT/_0514_ ), .A2(\CLINT/_0220_ ), .ZN(\CLINT/_0515_ ) );
OAI21_X1 \CLINT/_1240_ ( .A(\CLINT/_0467_ ), .B1(\CLINT/_0514_ ), .B2(\CLINT/_0220_ ), .ZN(\CLINT/_0516_ ) );
NOR2_X1 \CLINT/_1241_ ( .A1(\CLINT/_0515_ ), .A2(\CLINT/_0516_ ), .ZN(\CLINT/_0088_ ) );
AND3_X1 \CLINT/_1242_ ( .A1(\CLINT/_0514_ ), .A2(\CLINT/_0220_ ), .A3(\CLINT/_0221_ ), .ZN(\CLINT/_0517_ ) );
AOI21_X1 \CLINT/_1243_ ( .A(\CLINT/_0221_ ), .B1(\CLINT/_0514_ ), .B2(\CLINT/_0220_ ), .ZN(\CLINT/_0518_ ) );
NOR3_X1 \CLINT/_1244_ ( .A1(\CLINT/_0517_ ), .A2(\CLINT/_0518_ ), .A3(fanout_net_7 ), .ZN(\CLINT/_0089_ ) );
AND2_X1 \CLINT/_1245_ ( .A1(\CLINT/_0517_ ), .A2(\CLINT/_0222_ ), .ZN(\CLINT/_0519_ ) );
OAI21_X1 \CLINT/_1246_ ( .A(\CLINT/_0467_ ), .B1(\CLINT/_0517_ ), .B2(\CLINT/_0222_ ), .ZN(\CLINT/_0520_ ) );
NOR2_X1 \CLINT/_1247_ ( .A1(\CLINT/_0519_ ), .A2(\CLINT/_0520_ ), .ZN(\CLINT/_0090_ ) );
AOI21_X1 \CLINT/_1248_ ( .A(\CLINT/_0223_ ), .B1(\CLINT/_0517_ ), .B2(\CLINT/_0222_ ), .ZN(\CLINT/_0521_ ) );
AND2_X1 \CLINT/_1249_ ( .A1(\CLINT/_0474_ ), .A2(\CLINT/_0500_ ), .ZN(\CLINT/_0522_ ) );
AND4_X1 \CLINT/_1250_ ( .A1(\CLINT/_0220_ ), .A2(\CLINT/_0221_ ), .A3(\CLINT/_0222_ ), .A4(\CLINT/_0223_ ), .ZN(\CLINT/_0523_ ) );
AND3_X1 \CLINT/_1251_ ( .A1(\CLINT/_0523_ ), .A2(\CLINT/_0506_ ), .A3(\CLINT/_0512_ ), .ZN(\CLINT/_0524_ ) );
AND2_X1 \CLINT/_1252_ ( .A1(\CLINT/_0522_ ), .A2(\CLINT/_0524_ ), .ZN(\CLINT/_0525_ ) );
NOR3_X1 \CLINT/_1253_ ( .A1(\CLINT/_0521_ ), .A2(fanout_net_7 ), .A3(\CLINT/_0525_ ), .ZN(\CLINT/_0091_ ) );
AND3_X4 \CLINT/_1254_ ( .A1(\CLINT/_0452_ ), .A2(\CLINT/_0500_ ), .A3(\CLINT/_0524_ ), .ZN(\CLINT/_0526_ ) );
AND2_X1 \CLINT/_1255_ ( .A1(\CLINT/_0526_ ), .A2(\CLINT/_0224_ ), .ZN(\CLINT/_0527_ ) );
OAI21_X1 \CLINT/_1256_ ( .A(\CLINT/_0467_ ), .B1(\CLINT/_0526_ ), .B2(\CLINT/_0224_ ), .ZN(\CLINT/_0528_ ) );
NOR2_X1 \CLINT/_1257_ ( .A1(\CLINT/_0527_ ), .A2(\CLINT/_0528_ ), .ZN(\CLINT/_0092_ ) );
AND3_X1 \CLINT/_1258_ ( .A1(\CLINT/_0526_ ), .A2(\CLINT/_0224_ ), .A3(\CLINT/_0225_ ), .ZN(\CLINT/_0529_ ) );
AOI21_X1 \CLINT/_1259_ ( .A(\CLINT/_0225_ ), .B1(\CLINT/_0526_ ), .B2(\CLINT/_0224_ ), .ZN(\CLINT/_0530_ ) );
NOR3_X1 \CLINT/_1260_ ( .A1(\CLINT/_0529_ ), .A2(\CLINT/_0530_ ), .A3(fanout_net_7 ), .ZN(\CLINT/_0093_ ) );
AND2_X1 \CLINT/_1261_ ( .A1(\CLINT/_0529_ ), .A2(\CLINT/_0226_ ), .ZN(\CLINT/_0531_ ) );
OAI21_X1 \CLINT/_1262_ ( .A(\CLINT/_0467_ ), .B1(\CLINT/_0529_ ), .B2(\CLINT/_0226_ ), .ZN(\CLINT/_0532_ ) );
NOR2_X1 \CLINT/_1263_ ( .A1(\CLINT/_0531_ ), .A2(\CLINT/_0532_ ), .ZN(\CLINT/_0094_ ) );
AND3_X1 \CLINT/_1264_ ( .A1(\CLINT/_0529_ ), .A2(\CLINT/_0226_ ), .A3(\CLINT/_0227_ ), .ZN(\CLINT/_0533_ ) );
AOI21_X1 \CLINT/_1265_ ( .A(\CLINT/_0227_ ), .B1(\CLINT/_0529_ ), .B2(\CLINT/_0226_ ), .ZN(\CLINT/_0534_ ) );
NOR3_X1 \CLINT/_1266_ ( .A1(\CLINT/_0533_ ), .A2(\CLINT/_0534_ ), .A3(\CLINT/_0577_ ), .ZN(\CLINT/_0095_ ) );
AND2_X1 \CLINT/_1267_ ( .A1(\CLINT/_0224_ ), .A2(\CLINT/_0225_ ), .ZN(\CLINT/_0535_ ) );
AND2_X1 \CLINT/_1268_ ( .A1(\CLINT/_0226_ ), .A2(\CLINT/_0227_ ), .ZN(\CLINT/_0536_ ) );
AND3_X4 \CLINT/_1269_ ( .A1(\CLINT/_0526_ ), .A2(\CLINT/_0535_ ), .A3(\CLINT/_0536_ ), .ZN(\CLINT/_0537_ ) );
AND2_X1 \CLINT/_1270_ ( .A1(\CLINT/_0537_ ), .A2(\CLINT/_0229_ ), .ZN(\CLINT/_0538_ ) );
OAI21_X1 \CLINT/_1271_ ( .A(\CLINT/_0467_ ), .B1(\CLINT/_0537_ ), .B2(\CLINT/_0229_ ), .ZN(\CLINT/_0539_ ) );
NOR2_X1 \CLINT/_1272_ ( .A1(\CLINT/_0538_ ), .A2(\CLINT/_0539_ ), .ZN(\CLINT/_0096_ ) );
AND3_X4 \CLINT/_1273_ ( .A1(\CLINT/_0537_ ), .A2(\CLINT/_0229_ ), .A3(\CLINT/_0230_ ), .ZN(\CLINT/_0540_ ) );
AOI21_X1 \CLINT/_1274_ ( .A(\CLINT/_0230_ ), .B1(\CLINT/_0537_ ), .B2(\CLINT/_0229_ ), .ZN(\CLINT/_0541_ ) );
NOR3_X1 \CLINT/_1275_ ( .A1(\CLINT/_0540_ ), .A2(\CLINT/_0541_ ), .A3(\CLINT/_0577_ ), .ZN(\CLINT/_0097_ ) );
AND3_X4 \CLINT/_1276_ ( .A1(\CLINT/_0537_ ), .A2(\CLINT/_0229_ ), .A3(\CLINT/_0230_ ), .ZN(\CLINT/_0542_ ) );
AND2_X1 \CLINT/_1277_ ( .A1(\CLINT/_0542_ ), .A2(\CLINT/_0231_ ), .ZN(\CLINT/_0543_ ) );
OAI21_X1 \CLINT/_1278_ ( .A(\CLINT/_0467_ ), .B1(\CLINT/_0540_ ), .B2(\CLINT/_0231_ ), .ZN(\CLINT/_0544_ ) );
NOR2_X1 \CLINT/_1279_ ( .A1(\CLINT/_0543_ ), .A2(\CLINT/_0544_ ), .ZN(\CLINT/_0098_ ) );
AND3_X2 \CLINT/_1280_ ( .A1(\CLINT/_0542_ ), .A2(\CLINT/_0231_ ), .A3(\CLINT/_0232_ ), .ZN(\CLINT/_0545_ ) );
AOI21_X2 \CLINT/_1281_ ( .A(\CLINT/_0232_ ), .B1(\CLINT/_0542_ ), .B2(\CLINT/_0231_ ), .ZN(\CLINT/_0546_ ) );
NOR3_X1 \CLINT/_1282_ ( .A1(\CLINT/_0545_ ), .A2(\CLINT/_0546_ ), .A3(\CLINT/_0577_ ), .ZN(\CLINT/_0099_ ) );
DFF_X1 \CLINT/_1283_ ( .D(\CLINT/_0741_ ), .CK(clock ), .Q(\CLINT/state [0] ), .QN(\CLINT/_0740_ ) );
DFF_X1 \CLINT/_1284_ ( .D(\CLINT/_0742_ ), .CK(clock ), .Q(\CLINT/state [1] ), .QN(\CLINT/_0739_ ) );
DFF_X1 \CLINT/_1285_ ( .D(\CLINT/_0743_ ), .CK(clock ), .Q(\CLINT/readAddr [2] ), .QN(\CLINT/_0738_ ) );
DFF_X1 \CLINT/_1286_ ( .D(\CLINT/_0744_ ), .CK(clock ), .Q(\CLINT/readAddr [3] ), .QN(\CLINT/_0737_ ) );
DFF_X1 \CLINT/_1287_ ( .D(\CLINT/_0745_ ), .CK(clock ), .Q(\CLINT/readAddr [4] ), .QN(\CLINT/_0736_ ) );
DFF_X1 \CLINT/_1288_ ( .D(\CLINT/_0746_ ), .CK(clock ), .Q(\CLINT/readAddr [5] ), .QN(\CLINT/_0735_ ) );
DFF_X1 \CLINT/_1289_ ( .D(\CLINT/_0747_ ), .CK(clock ), .Q(\CLINT/readAddr [6] ), .QN(\CLINT/_0734_ ) );
DFF_X1 \CLINT/_1290_ ( .D(\CLINT/_0748_ ), .CK(clock ), .Q(\CLINT/readAddr [7] ), .QN(\CLINT/_0733_ ) );
DFF_X1 \CLINT/_1291_ ( .D(\CLINT/_0749_ ), .CK(clock ), .Q(\CLINT/readAddr [8] ), .QN(\CLINT/_0732_ ) );
DFF_X1 \CLINT/_1292_ ( .D(\CLINT/_0750_ ), .CK(clock ), .Q(\CLINT/readAddr [9] ), .QN(\CLINT/_0731_ ) );
DFF_X1 \CLINT/_1293_ ( .D(\CLINT/_0751_ ), .CK(clock ), .Q(\CLINT/readAddr [10] ), .QN(\CLINT/_0730_ ) );
DFF_X1 \CLINT/_1294_ ( .D(\CLINT/_0752_ ), .CK(clock ), .Q(\CLINT/readAddr [11] ), .QN(\CLINT/_0729_ ) );
DFF_X1 \CLINT/_1295_ ( .D(\CLINT/_0753_ ), .CK(clock ), .Q(\CLINT/readAddr [12] ), .QN(\CLINT/_0728_ ) );
DFF_X1 \CLINT/_1296_ ( .D(\CLINT/_0754_ ), .CK(clock ), .Q(\CLINT/readAddr [13] ), .QN(\CLINT/_0727_ ) );
DFF_X1 \CLINT/_1297_ ( .D(\CLINT/_0755_ ), .CK(clock ), .Q(\CLINT/readAddr [14] ), .QN(\CLINT/_0726_ ) );
DFF_X1 \CLINT/_1298_ ( .D(\CLINT/_0756_ ), .CK(clock ), .Q(\CLINT/readAddr [15] ), .QN(\CLINT/_0725_ ) );
DFF_X1 \CLINT/_1299_ ( .D(\CLINT/_0757_ ), .CK(clock ), .Q(\CLINT/readAddr [16] ), .QN(\CLINT/_0724_ ) );
DFF_X1 \CLINT/_1300_ ( .D(\CLINT/_0758_ ), .CK(clock ), .Q(\CLINT/readAddr [17] ), .QN(\CLINT/_0723_ ) );
DFF_X1 \CLINT/_1301_ ( .D(\CLINT/_0759_ ), .CK(clock ), .Q(\CLINT/readAddr [18] ), .QN(\CLINT/_0722_ ) );
DFF_X1 \CLINT/_1302_ ( .D(\CLINT/_0760_ ), .CK(clock ), .Q(\CLINT/readAddr [19] ), .QN(\CLINT/_0721_ ) );
DFF_X1 \CLINT/_1303_ ( .D(\CLINT/_0761_ ), .CK(clock ), .Q(\CLINT/readAddr [20] ), .QN(\CLINT/_0720_ ) );
DFF_X1 \CLINT/_1304_ ( .D(\CLINT/_0762_ ), .CK(clock ), .Q(\CLINT/readAddr [21] ), .QN(\CLINT/_0719_ ) );
DFF_X1 \CLINT/_1305_ ( .D(\CLINT/_0763_ ), .CK(clock ), .Q(\CLINT/readAddr [22] ), .QN(\CLINT/_0718_ ) );
DFF_X1 \CLINT/_1306_ ( .D(\CLINT/_0764_ ), .CK(clock ), .Q(\CLINT/readAddr [23] ), .QN(\CLINT/_0717_ ) );
DFF_X1 \CLINT/_1307_ ( .D(\CLINT/_0765_ ), .CK(clock ), .Q(\CLINT/readAddr [24] ), .QN(\CLINT/_0716_ ) );
DFF_X1 \CLINT/_1308_ ( .D(\CLINT/_0766_ ), .CK(clock ), .Q(\CLINT/readAddr [25] ), .QN(\CLINT/_0715_ ) );
DFF_X1 \CLINT/_1309_ ( .D(\CLINT/_0767_ ), .CK(clock ), .Q(\CLINT/readAddr [26] ), .QN(\CLINT/_0714_ ) );
DFF_X1 \CLINT/_1310_ ( .D(\CLINT/_0768_ ), .CK(clock ), .Q(\CLINT/readAddr [27] ), .QN(\CLINT/_0713_ ) );
DFF_X1 \CLINT/_1311_ ( .D(\CLINT/_0769_ ), .CK(clock ), .Q(\CLINT/readAddr [28] ), .QN(\CLINT/_0712_ ) );
DFF_X1 \CLINT/_1312_ ( .D(\CLINT/_0770_ ), .CK(clock ), .Q(\CLINT/readAddr [29] ), .QN(\CLINT/_0711_ ) );
DFF_X1 \CLINT/_1313_ ( .D(\CLINT/_0771_ ), .CK(clock ), .Q(\CLINT/readAddr [30] ), .QN(\CLINT/_0710_ ) );
DFF_X1 \CLINT/_1314_ ( .D(\CLINT/_0772_ ), .CK(clock ), .Q(\CLINT/readAddr [31] ), .QN(\CLINT/_0709_ ) );
DFF_X1 \CLINT/_1315_ ( .D(\CLINT/_0773_ ), .CK(clock ), .Q(\CLINT/state [2] ), .QN(\CLINT/_0000_ ) );
DFF_X1 \CLINT/_1316_ ( .D(\CLINT/_0774_ ), .CK(clock ), .Q(\CLINT/mtime [0] ), .QN(\CLINT/_0581_ ) );
DFF_X1 \CLINT/_1317_ ( .D(\CLINT/_0775_ ), .CK(clock ), .Q(\CLINT/mtime [1] ), .QN(\CLINT/_0708_ ) );
DFF_X1 \CLINT/_1318_ ( .D(\CLINT/_0776_ ), .CK(clock ), .Q(\CLINT/mtime [2] ), .QN(\CLINT/_0707_ ) );
DFF_X1 \CLINT/_1319_ ( .D(\CLINT/_0777_ ), .CK(clock ), .Q(\CLINT/mtime [3] ), .QN(\CLINT/_0706_ ) );
DFF_X1 \CLINT/_1320_ ( .D(\CLINT/_0778_ ), .CK(clock ), .Q(\CLINT/mtime [4] ), .QN(\CLINT/_0705_ ) );
DFF_X1 \CLINT/_1321_ ( .D(\CLINT/_0779_ ), .CK(clock ), .Q(\CLINT/mtime [5] ), .QN(\CLINT/_0704_ ) );
DFF_X1 \CLINT/_1322_ ( .D(\CLINT/_0780_ ), .CK(clock ), .Q(\CLINT/mtime [6] ), .QN(\CLINT/_0703_ ) );
DFF_X1 \CLINT/_1323_ ( .D(\CLINT/_0781_ ), .CK(clock ), .Q(\CLINT/mtime [7] ), .QN(\CLINT/_0702_ ) );
DFF_X1 \CLINT/_1324_ ( .D(\CLINT/_0782_ ), .CK(clock ), .Q(\CLINT/mtime [8] ), .QN(\CLINT/_0701_ ) );
DFF_X1 \CLINT/_1325_ ( .D(\CLINT/_0783_ ), .CK(clock ), .Q(\CLINT/mtime [9] ), .QN(\CLINT/_0700_ ) );
DFF_X1 \CLINT/_1326_ ( .D(\CLINT/_0784_ ), .CK(clock ), .Q(\CLINT/mtime [10] ), .QN(\CLINT/_0699_ ) );
DFF_X1 \CLINT/_1327_ ( .D(\CLINT/_0785_ ), .CK(clock ), .Q(\CLINT/mtime [11] ), .QN(\CLINT/_0698_ ) );
DFF_X1 \CLINT/_1328_ ( .D(\CLINT/_0786_ ), .CK(clock ), .Q(\CLINT/mtime [12] ), .QN(\CLINT/_0697_ ) );
DFF_X1 \CLINT/_1329_ ( .D(\CLINT/_0787_ ), .CK(clock ), .Q(\CLINT/mtime [13] ), .QN(\CLINT/_0696_ ) );
DFF_X1 \CLINT/_1330_ ( .D(\CLINT/_0788_ ), .CK(clock ), .Q(\CLINT/mtime [14] ), .QN(\CLINT/_0695_ ) );
DFF_X1 \CLINT/_1331_ ( .D(\CLINT/_0789_ ), .CK(clock ), .Q(\CLINT/mtime [15] ), .QN(\CLINT/_0694_ ) );
DFF_X1 \CLINT/_1332_ ( .D(\CLINT/_0790_ ), .CK(clock ), .Q(\CLINT/mtime [16] ), .QN(\CLINT/_0693_ ) );
DFF_X1 \CLINT/_1333_ ( .D(\CLINT/_0791_ ), .CK(clock ), .Q(\CLINT/mtime [17] ), .QN(\CLINT/_0692_ ) );
DFF_X1 \CLINT/_1334_ ( .D(\CLINT/_0792_ ), .CK(clock ), .Q(\CLINT/mtime [18] ), .QN(\CLINT/_0691_ ) );
DFF_X1 \CLINT/_1335_ ( .D(\CLINT/_0793_ ), .CK(clock ), .Q(\CLINT/mtime [19] ), .QN(\CLINT/_0690_ ) );
DFF_X1 \CLINT/_1336_ ( .D(\CLINT/_0794_ ), .CK(clock ), .Q(\CLINT/mtime [20] ), .QN(\CLINT/_0689_ ) );
DFF_X1 \CLINT/_1337_ ( .D(\CLINT/_0795_ ), .CK(clock ), .Q(\CLINT/mtime [21] ), .QN(\CLINT/_0688_ ) );
DFF_X1 \CLINT/_1338_ ( .D(\CLINT/_0796_ ), .CK(clock ), .Q(\CLINT/mtime [22] ), .QN(\CLINT/_0687_ ) );
DFF_X1 \CLINT/_1339_ ( .D(\CLINT/_0797_ ), .CK(clock ), .Q(\CLINT/mtime [23] ), .QN(\CLINT/_0686_ ) );
DFF_X1 \CLINT/_1340_ ( .D(\CLINT/_0798_ ), .CK(clock ), .Q(\CLINT/mtime [24] ), .QN(\CLINT/_0685_ ) );
DFF_X1 \CLINT/_1341_ ( .D(\CLINT/_0799_ ), .CK(clock ), .Q(\CLINT/mtime [25] ), .QN(\CLINT/_0684_ ) );
DFF_X1 \CLINT/_1342_ ( .D(\CLINT/_0800_ ), .CK(clock ), .Q(\CLINT/mtime [26] ), .QN(\CLINT/_0683_ ) );
DFF_X1 \CLINT/_1343_ ( .D(\CLINT/_0801_ ), .CK(clock ), .Q(\CLINT/mtime [27] ), .QN(\CLINT/_0682_ ) );
DFF_X1 \CLINT/_1344_ ( .D(\CLINT/_0802_ ), .CK(clock ), .Q(\CLINT/mtime [28] ), .QN(\CLINT/_0681_ ) );
DFF_X1 \CLINT/_1345_ ( .D(\CLINT/_0803_ ), .CK(clock ), .Q(\CLINT/mtime [29] ), .QN(\CLINT/_0680_ ) );
DFF_X1 \CLINT/_1346_ ( .D(\CLINT/_0804_ ), .CK(clock ), .Q(\CLINT/mtime [30] ), .QN(\CLINT/_0679_ ) );
DFF_X1 \CLINT/_1347_ ( .D(\CLINT/_0805_ ), .CK(clock ), .Q(\CLINT/mtime [31] ), .QN(\CLINT/_0678_ ) );
DFF_X1 \CLINT/_1348_ ( .D(\CLINT/_0806_ ), .CK(clock ), .Q(\CLINT/mtime [32] ), .QN(\CLINT/_0677_ ) );
DFF_X1 \CLINT/_1349_ ( .D(\CLINT/_0807_ ), .CK(clock ), .Q(\CLINT/mtime [33] ), .QN(\CLINT/_0676_ ) );
DFF_X1 \CLINT/_1350_ ( .D(\CLINT/_0808_ ), .CK(clock ), .Q(\CLINT/mtime [34] ), .QN(\CLINT/_0675_ ) );
DFF_X1 \CLINT/_1351_ ( .D(\CLINT/_0809_ ), .CK(clock ), .Q(\CLINT/mtime [35] ), .QN(\CLINT/_0674_ ) );
DFF_X1 \CLINT/_1352_ ( .D(\CLINT/_0810_ ), .CK(clock ), .Q(\CLINT/mtime [36] ), .QN(\CLINT/_0673_ ) );
DFF_X1 \CLINT/_1353_ ( .D(\CLINT/_0811_ ), .CK(clock ), .Q(\CLINT/mtime [37] ), .QN(\CLINT/_0672_ ) );
DFF_X1 \CLINT/_1354_ ( .D(\CLINT/_0812_ ), .CK(clock ), .Q(\CLINT/mtime [38] ), .QN(\CLINT/_0671_ ) );
DFF_X1 \CLINT/_1355_ ( .D(\CLINT/_0813_ ), .CK(clock ), .Q(\CLINT/mtime [39] ), .QN(\CLINT/_0670_ ) );
DFF_X1 \CLINT/_1356_ ( .D(\CLINT/_0814_ ), .CK(clock ), .Q(\CLINT/mtime [40] ), .QN(\CLINT/_0669_ ) );
DFF_X1 \CLINT/_1357_ ( .D(\CLINT/_0815_ ), .CK(clock ), .Q(\CLINT/mtime [41] ), .QN(\CLINT/_0668_ ) );
DFF_X1 \CLINT/_1358_ ( .D(\CLINT/_0816_ ), .CK(clock ), .Q(\CLINT/mtime [42] ), .QN(\CLINT/_0667_ ) );
DFF_X1 \CLINT/_1359_ ( .D(\CLINT/_0817_ ), .CK(clock ), .Q(\CLINT/mtime [43] ), .QN(\CLINT/_0666_ ) );
DFF_X1 \CLINT/_1360_ ( .D(\CLINT/_0818_ ), .CK(clock ), .Q(\CLINT/mtime [44] ), .QN(\CLINT/_0665_ ) );
DFF_X1 \CLINT/_1361_ ( .D(\CLINT/_0819_ ), .CK(clock ), .Q(\CLINT/mtime [45] ), .QN(\CLINT/_0664_ ) );
DFF_X1 \CLINT/_1362_ ( .D(\CLINT/_0820_ ), .CK(clock ), .Q(\CLINT/mtime [46] ), .QN(\CLINT/_0663_ ) );
DFF_X1 \CLINT/_1363_ ( .D(\CLINT/_0821_ ), .CK(clock ), .Q(\CLINT/mtime [47] ), .QN(\CLINT/_0662_ ) );
DFF_X1 \CLINT/_1364_ ( .D(\CLINT/_0822_ ), .CK(clock ), .Q(\CLINT/mtime [48] ), .QN(\CLINT/_0661_ ) );
DFF_X1 \CLINT/_1365_ ( .D(\CLINT/_0823_ ), .CK(clock ), .Q(\CLINT/mtime [49] ), .QN(\CLINT/_0660_ ) );
DFF_X1 \CLINT/_1366_ ( .D(\CLINT/_0824_ ), .CK(clock ), .Q(\CLINT/mtime [50] ), .QN(\CLINT/_0659_ ) );
DFF_X1 \CLINT/_1367_ ( .D(\CLINT/_0825_ ), .CK(clock ), .Q(\CLINT/mtime [51] ), .QN(\CLINT/_0658_ ) );
DFF_X1 \CLINT/_1368_ ( .D(\CLINT/_0826_ ), .CK(clock ), .Q(\CLINT/mtime [52] ), .QN(\CLINT/_0657_ ) );
DFF_X1 \CLINT/_1369_ ( .D(\CLINT/_0827_ ), .CK(clock ), .Q(\CLINT/mtime [53] ), .QN(\CLINT/_0656_ ) );
DFF_X1 \CLINT/_1370_ ( .D(\CLINT/_0828_ ), .CK(clock ), .Q(\CLINT/mtime [54] ), .QN(\CLINT/_0655_ ) );
DFF_X1 \CLINT/_1371_ ( .D(\CLINT/_0829_ ), .CK(clock ), .Q(\CLINT/mtime [55] ), .QN(\CLINT/_0654_ ) );
DFF_X1 \CLINT/_1372_ ( .D(\CLINT/_0830_ ), .CK(clock ), .Q(\CLINT/mtime [56] ), .QN(\CLINT/_0653_ ) );
DFF_X1 \CLINT/_1373_ ( .D(\CLINT/_0831_ ), .CK(clock ), .Q(\CLINT/mtime [57] ), .QN(\CLINT/_0652_ ) );
DFF_X1 \CLINT/_1374_ ( .D(\CLINT/_0832_ ), .CK(clock ), .Q(\CLINT/mtime [58] ), .QN(\CLINT/_0651_ ) );
DFF_X1 \CLINT/_1375_ ( .D(\CLINT/_0833_ ), .CK(clock ), .Q(\CLINT/mtime [59] ), .QN(\CLINT/_0650_ ) );
DFF_X1 \CLINT/_1376_ ( .D(\CLINT/_0834_ ), .CK(clock ), .Q(\CLINT/mtime [60] ), .QN(\CLINT/_0649_ ) );
DFF_X1 \CLINT/_1377_ ( .D(\CLINT/_0835_ ), .CK(clock ), .Q(\CLINT/mtime [61] ), .QN(\CLINT/_0648_ ) );
DFF_X1 \CLINT/_1378_ ( .D(\CLINT/_0836_ ), .CK(clock ), .Q(\CLINT/mtime [62] ), .QN(\CLINT/_0647_ ) );
DFF_X1 \CLINT/_1379_ ( .D(\CLINT/_0837_ ), .CK(clock ), .Q(\CLINT/mtime [63] ), .QN(\CLINT/_0646_ ) );
BUF_X1 \CLINT/_1380_ ( .A(\CLINT/mtime [1] ), .Z(\CLINT/_0592_ ) );
BUF_X1 \CLINT/_1381_ ( .A(\CLINT/mtime [2] ), .Z(\CLINT/_0603_ ) );
BUF_X1 \CLINT/_1382_ ( .A(\CLINT/mtime [3] ), .Z(\CLINT/_0614_ ) );
BUF_X1 \CLINT/_1383_ ( .A(\CLINT/mtime [4] ), .Z(\CLINT/_0625_ ) );
BUF_X1 \CLINT/_1384_ ( .A(\CLINT/mtime [5] ), .Z(\CLINT/_0636_ ) );
BUF_X1 \CLINT/_1385_ ( .A(\CLINT/mtime [6] ), .Z(\CLINT/_0641_ ) );
BUF_X1 \CLINT/_1386_ ( .A(\CLINT/mtime [7] ), .Z(\CLINT/_0642_ ) );
BUF_X1 \CLINT/_1387_ ( .A(\CLINT/mtime [8] ), .Z(\CLINT/_0643_ ) );
BUF_X1 \CLINT/_1388_ ( .A(\CLINT/mtime [9] ), .Z(\CLINT/_0644_ ) );
BUF_X1 \CLINT/_1389_ ( .A(\CLINT/mtime [10] ), .Z(\CLINT/_0582_ ) );
BUF_X1 \CLINT/_1390_ ( .A(\CLINT/mtime [11] ), .Z(\CLINT/_0583_ ) );
BUF_X1 \CLINT/_1391_ ( .A(\CLINT/mtime [12] ), .Z(\CLINT/_0584_ ) );
BUF_X1 \CLINT/_1392_ ( .A(\CLINT/mtime [13] ), .Z(\CLINT/_0585_ ) );
BUF_X1 \CLINT/_1393_ ( .A(\CLINT/mtime [14] ), .Z(\CLINT/_0586_ ) );
BUF_X1 \CLINT/_1394_ ( .A(\CLINT/mtime [15] ), .Z(\CLINT/_0587_ ) );
BUF_X1 \CLINT/_1395_ ( .A(\CLINT/mtime [16] ), .Z(\CLINT/_0588_ ) );
BUF_X1 \CLINT/_1396_ ( .A(\CLINT/mtime [17] ), .Z(\CLINT/_0589_ ) );
BUF_X1 \CLINT/_1397_ ( .A(\CLINT/mtime [18] ), .Z(\CLINT/_0590_ ) );
BUF_X1 \CLINT/_1398_ ( .A(\CLINT/mtime [19] ), .Z(\CLINT/_0591_ ) );
BUF_X1 \CLINT/_1399_ ( .A(\CLINT/mtime [20] ), .Z(\CLINT/_0593_ ) );
BUF_X1 \CLINT/_1400_ ( .A(\CLINT/mtime [21] ), .Z(\CLINT/_0594_ ) );
BUF_X1 \CLINT/_1401_ ( .A(\CLINT/mtime [22] ), .Z(\CLINT/_0595_ ) );
BUF_X1 \CLINT/_1402_ ( .A(\CLINT/mtime [23] ), .Z(\CLINT/_0596_ ) );
BUF_X1 \CLINT/_1403_ ( .A(\CLINT/mtime [24] ), .Z(\CLINT/_0597_ ) );
BUF_X1 \CLINT/_1404_ ( .A(\CLINT/mtime [25] ), .Z(\CLINT/_0598_ ) );
BUF_X1 \CLINT/_1405_ ( .A(\CLINT/mtime [26] ), .Z(\CLINT/_0599_ ) );
BUF_X1 \CLINT/_1406_ ( .A(\CLINT/mtime [27] ), .Z(\CLINT/_0600_ ) );
BUF_X1 \CLINT/_1407_ ( .A(\CLINT/mtime [28] ), .Z(\CLINT/_0601_ ) );
BUF_X1 \CLINT/_1408_ ( .A(\CLINT/mtime [29] ), .Z(\CLINT/_0602_ ) );
BUF_X1 \CLINT/_1409_ ( .A(\CLINT/mtime [30] ), .Z(\CLINT/_0604_ ) );
BUF_X1 \CLINT/_1410_ ( .A(\CLINT/mtime [31] ), .Z(\CLINT/_0605_ ) );
BUF_X1 \CLINT/_1411_ ( .A(\CLINT/mtime [32] ), .Z(\CLINT/_0606_ ) );
BUF_X1 \CLINT/_1412_ ( .A(\CLINT/mtime [33] ), .Z(\CLINT/_0607_ ) );
BUF_X1 \CLINT/_1413_ ( .A(\CLINT/mtime [34] ), .Z(\CLINT/_0608_ ) );
BUF_X1 \CLINT/_1414_ ( .A(\CLINT/mtime [35] ), .Z(\CLINT/_0609_ ) );
BUF_X1 \CLINT/_1415_ ( .A(\CLINT/mtime [36] ), .Z(\CLINT/_0610_ ) );
BUF_X1 \CLINT/_1416_ ( .A(\CLINT/mtime [37] ), .Z(\CLINT/_0611_ ) );
BUF_X1 \CLINT/_1417_ ( .A(\CLINT/mtime [38] ), .Z(\CLINT/_0612_ ) );
BUF_X1 \CLINT/_1418_ ( .A(\CLINT/mtime [39] ), .Z(\CLINT/_0613_ ) );
BUF_X1 \CLINT/_1419_ ( .A(\CLINT/mtime [40] ), .Z(\CLINT/_0615_ ) );
BUF_X1 \CLINT/_1420_ ( .A(\CLINT/mtime [41] ), .Z(\CLINT/_0616_ ) );
BUF_X1 \CLINT/_1421_ ( .A(\CLINT/mtime [42] ), .Z(\CLINT/_0617_ ) );
BUF_X1 \CLINT/_1422_ ( .A(\CLINT/mtime [43] ), .Z(\CLINT/_0618_ ) );
BUF_X1 \CLINT/_1423_ ( .A(\CLINT/mtime [44] ), .Z(\CLINT/_0619_ ) );
BUF_X1 \CLINT/_1424_ ( .A(\CLINT/mtime [45] ), .Z(\CLINT/_0620_ ) );
BUF_X1 \CLINT/_1425_ ( .A(\CLINT/mtime [46] ), .Z(\CLINT/_0621_ ) );
BUF_X1 \CLINT/_1426_ ( .A(\CLINT/mtime [47] ), .Z(\CLINT/_0622_ ) );
BUF_X1 \CLINT/_1427_ ( .A(\CLINT/mtime [48] ), .Z(\CLINT/_0623_ ) );
BUF_X1 \CLINT/_1428_ ( .A(\CLINT/mtime [49] ), .Z(\CLINT/_0624_ ) );
BUF_X1 \CLINT/_1429_ ( .A(\CLINT/mtime [50] ), .Z(\CLINT/_0626_ ) );
BUF_X1 \CLINT/_1430_ ( .A(\CLINT/mtime [51] ), .Z(\CLINT/_0627_ ) );
BUF_X1 \CLINT/_1431_ ( .A(\CLINT/mtime [52] ), .Z(\CLINT/_0628_ ) );
BUF_X1 \CLINT/_1432_ ( .A(\CLINT/mtime [53] ), .Z(\CLINT/_0629_ ) );
BUF_X1 \CLINT/_1433_ ( .A(\CLINT/mtime [54] ), .Z(\CLINT/_0630_ ) );
BUF_X1 \CLINT/_1434_ ( .A(\CLINT/mtime [55] ), .Z(\CLINT/_0631_ ) );
BUF_X1 \CLINT/_1435_ ( .A(\CLINT/mtime [56] ), .Z(\CLINT/_0632_ ) );
BUF_X1 \CLINT/_1436_ ( .A(\CLINT/mtime [57] ), .Z(\CLINT/_0633_ ) );
BUF_X1 \CLINT/_1437_ ( .A(\CLINT/mtime [58] ), .Z(\CLINT/_0634_ ) );
BUF_X1 \CLINT/_1438_ ( .A(\CLINT/mtime [59] ), .Z(\CLINT/_0635_ ) );
BUF_X1 \CLINT/_1439_ ( .A(\CLINT/mtime [60] ), .Z(\CLINT/_0637_ ) );
BUF_X1 \CLINT/_1440_ ( .A(\CLINT/mtime [61] ), .Z(\CLINT/_0638_ ) );
BUF_X1 \CLINT/_1441_ ( .A(\CLINT/mtime [62] ), .Z(\CLINT/_0639_ ) );
BUF_X1 \CLINT/_1442_ ( .A(\CLINT/mtime [63] ), .Z(\CLINT/_0640_ ) );
BUF_X1 \CLINT/_1443_ ( .A(\CLINT/_0581_ ), .Z(\CLINT/_0645_ ) );
BUF_X1 \CLINT/_1444_ ( .A(_CLINT_io_bvalid ), .Z(\_CLINT_io_bresp [0] ) );
BUF_X1 \CLINT/_1445_ ( .A(_CLINT_io_bvalid ), .Z(\_CLINT_io_bresp [1] ) );
BUF_X1 \CLINT/_1446_ ( .A(\_CLINT_io_rresp [1] ), .Z(\_CLINT_io_rresp [0] ) );
BUF_X1 \CLINT/_1447_ ( .A(\CLINT/state [0] ), .Z(\CLINT/_0578_ ) );
BUF_X1 \CLINT/_1448_ ( .A(\CLINT/state [1] ), .Z(\CLINT/_0579_ ) );
BUF_X1 \CLINT/_1449_ ( .A(\CLINT/state [2] ), .Z(\CLINT/_0580_ ) );
BUF_X1 \CLINT/_1450_ ( .A(\CLINT/_0170_ ), .Z(_CLINT_io_rvalid ) );
BUF_X1 \CLINT/_1451_ ( .A(reset ), .Z(\CLINT/_0577_ ) );
BUF_X1 \CLINT/_1452_ ( .A(\CLINT/_0000_ ), .Z(\CLINT/_0001_ ) );
BUF_X1 \CLINT/_1453_ ( .A(\CLINT/_0135_ ), .Z(_CLINT_io_bvalid ) );
BUF_X1 \CLINT/_1454_ ( .A(\CLINT/readAddr [2] ), .Z(\CLINT/_0567_ ) );
BUF_X1 \CLINT/_1455_ ( .A(\CLINT/readAddr [3] ), .Z(\CLINT/_0570_ ) );
BUF_X1 \CLINT/_1456_ ( .A(\CLINT/readAddr [5] ), .Z(\CLINT/_0572_ ) );
BUF_X1 \CLINT/_1457_ ( .A(\CLINT/readAddr [4] ), .Z(\CLINT/_0571_ ) );
BUF_X1 \CLINT/_1458_ ( .A(\CLINT/readAddr [7] ), .Z(\CLINT/_0574_ ) );
BUF_X1 \CLINT/_1459_ ( .A(\CLINT/readAddr [6] ), .Z(\CLINT/_0573_ ) );
BUF_X1 \CLINT/_1460_ ( .A(\CLINT/readAddr [9] ), .Z(\CLINT/_0576_ ) );
BUF_X1 \CLINT/_1461_ ( .A(\CLINT/readAddr [8] ), .Z(\CLINT/_0575_ ) );
BUF_X1 \CLINT/_1462_ ( .A(\CLINT/readAddr [11] ), .Z(\CLINT/_0548_ ) );
BUF_X1 \CLINT/_1463_ ( .A(\CLINT/readAddr [10] ), .Z(\CLINT/_0547_ ) );
BUF_X1 \CLINT/_1464_ ( .A(\CLINT/readAddr [13] ), .Z(\CLINT/_0550_ ) );
BUF_X1 \CLINT/_1465_ ( .A(\CLINT/readAddr [12] ), .Z(\CLINT/_0549_ ) );
BUF_X1 \CLINT/_1466_ ( .A(\CLINT/readAddr [15] ), .Z(\CLINT/_0552_ ) );
BUF_X1 \CLINT/_1467_ ( .A(\CLINT/readAddr [14] ), .Z(\CLINT/_0551_ ) );
BUF_X1 \CLINT/_1468_ ( .A(\CLINT/readAddr [17] ), .Z(\CLINT/_0554_ ) );
BUF_X1 \CLINT/_1469_ ( .A(\CLINT/readAddr [16] ), .Z(\CLINT/_0553_ ) );
BUF_X1 \CLINT/_1470_ ( .A(\CLINT/readAddr [19] ), .Z(\CLINT/_0556_ ) );
BUF_X1 \CLINT/_1471_ ( .A(\CLINT/readAddr [18] ), .Z(\CLINT/_0555_ ) );
BUF_X1 \CLINT/_1472_ ( .A(\CLINT/readAddr [21] ), .Z(\CLINT/_0558_ ) );
BUF_X1 \CLINT/_1473_ ( .A(\CLINT/readAddr [20] ), .Z(\CLINT/_0557_ ) );
BUF_X1 \CLINT/_1474_ ( .A(\CLINT/readAddr [23] ), .Z(\CLINT/_0560_ ) );
BUF_X1 \CLINT/_1475_ ( .A(\CLINT/readAddr [22] ), .Z(\CLINT/_0559_ ) );
BUF_X1 \CLINT/_1476_ ( .A(\CLINT/readAddr [24] ), .Z(\CLINT/_0561_ ) );
BUF_X1 \CLINT/_1477_ ( .A(\CLINT/readAddr [25] ), .Z(\CLINT/_0562_ ) );
BUF_X1 \CLINT/_1478_ ( .A(\CLINT/readAddr [27] ), .Z(\CLINT/_0564_ ) );
BUF_X1 \CLINT/_1479_ ( .A(\CLINT/readAddr [26] ), .Z(\CLINT/_0563_ ) );
BUF_X1 \CLINT/_1480_ ( .A(\CLINT/readAddr [29] ), .Z(\CLINT/_0566_ ) );
BUF_X1 \CLINT/_1481_ ( .A(\CLINT/readAddr [28] ), .Z(\CLINT/_0565_ ) );
BUF_X1 \CLINT/_1482_ ( .A(\CLINT/readAddr [31] ), .Z(\CLINT/_0569_ ) );
BUF_X1 \CLINT/_1483_ ( .A(\CLINT/readAddr [30] ), .Z(\CLINT/_0568_ ) );
BUF_X1 \CLINT/_1484_ ( .A(\CLINT/mtime [32] ), .Z(\CLINT/_0198_ ) );
BUF_X1 \CLINT/_1485_ ( .A(\CLINT/mtime [0] ), .Z(\CLINT/_0173_ ) );
BUF_X1 \CLINT/_1486_ ( .A(\CLINT/_0136_ ), .Z(\_CLINT_io_rdata [0] ) );
BUF_X1 \CLINT/_1487_ ( .A(\CLINT/mtime [33] ), .Z(\CLINT/_0199_ ) );
BUF_X1 \CLINT/_1488_ ( .A(\CLINT/mtime [1] ), .Z(\CLINT/_0184_ ) );
BUF_X1 \CLINT/_1489_ ( .A(\CLINT/_0147_ ), .Z(\_CLINT_io_rdata [1] ) );
BUF_X1 \CLINT/_1490_ ( .A(\CLINT/mtime [34] ), .Z(\CLINT/_0200_ ) );
BUF_X1 \CLINT/_1491_ ( .A(\CLINT/mtime [2] ), .Z(\CLINT/_0195_ ) );
BUF_X1 \CLINT/_1492_ ( .A(\CLINT/_0158_ ), .Z(\_CLINT_io_rdata [2] ) );
BUF_X1 \CLINT/_1493_ ( .A(\CLINT/mtime [35] ), .Z(\CLINT/_0201_ ) );
BUF_X1 \CLINT/_1494_ ( .A(\CLINT/mtime [3] ), .Z(\CLINT/_0206_ ) );
BUF_X1 \CLINT/_1495_ ( .A(\CLINT/_0161_ ), .Z(\_CLINT_io_rdata [3] ) );
BUF_X1 \CLINT/_1496_ ( .A(\CLINT/mtime [36] ), .Z(\CLINT/_0202_ ) );
BUF_X1 \CLINT/_1497_ ( .A(\CLINT/mtime [4] ), .Z(\CLINT/_0217_ ) );
BUF_X1 \CLINT/_1498_ ( .A(\CLINT/_0162_ ), .Z(\_CLINT_io_rdata [4] ) );
BUF_X1 \CLINT/_1499_ ( .A(\CLINT/mtime [37] ), .Z(\CLINT/_0203_ ) );
BUF_X1 \CLINT/_1500_ ( .A(\CLINT/mtime [5] ), .Z(\CLINT/_0228_ ) );
BUF_X1 \CLINT/_1501_ ( .A(\CLINT/_0163_ ), .Z(\_CLINT_io_rdata [5] ) );
BUF_X1 \CLINT/_1502_ ( .A(\CLINT/mtime [38] ), .Z(\CLINT/_0204_ ) );
BUF_X1 \CLINT/_1503_ ( .A(\CLINT/mtime [6] ), .Z(\CLINT/_0233_ ) );
BUF_X1 \CLINT/_1504_ ( .A(\CLINT/_0164_ ), .Z(\_CLINT_io_rdata [6] ) );
BUF_X1 \CLINT/_1505_ ( .A(\CLINT/mtime [39] ), .Z(\CLINT/_0205_ ) );
BUF_X1 \CLINT/_1506_ ( .A(\CLINT/mtime [7] ), .Z(\CLINT/_0234_ ) );
BUF_X1 \CLINT/_1507_ ( .A(\CLINT/_0165_ ), .Z(\_CLINT_io_rdata [7] ) );
BUF_X1 \CLINT/_1508_ ( .A(\CLINT/mtime [40] ), .Z(\CLINT/_0207_ ) );
BUF_X1 \CLINT/_1509_ ( .A(\CLINT/mtime [8] ), .Z(\CLINT/_0235_ ) );
BUF_X1 \CLINT/_1510_ ( .A(\CLINT/_0166_ ), .Z(\_CLINT_io_rdata [8] ) );
BUF_X1 \CLINT/_1511_ ( .A(\CLINT/mtime [41] ), .Z(\CLINT/_0208_ ) );
BUF_X1 \CLINT/_1512_ ( .A(\CLINT/mtime [9] ), .Z(\CLINT/_0236_ ) );
BUF_X1 \CLINT/_1513_ ( .A(\CLINT/_0167_ ), .Z(\_CLINT_io_rdata [9] ) );
BUF_X1 \CLINT/_1514_ ( .A(\CLINT/mtime [42] ), .Z(\CLINT/_0209_ ) );
BUF_X1 \CLINT/_1515_ ( .A(\CLINT/mtime [10] ), .Z(\CLINT/_0174_ ) );
BUF_X1 \CLINT/_1516_ ( .A(\CLINT/_0137_ ), .Z(\_CLINT_io_rdata [10] ) );
BUF_X1 \CLINT/_1517_ ( .A(\CLINT/mtime [43] ), .Z(\CLINT/_0210_ ) );
BUF_X1 \CLINT/_1518_ ( .A(\CLINT/mtime [11] ), .Z(\CLINT/_0175_ ) );
BUF_X1 \CLINT/_1519_ ( .A(\CLINT/_0138_ ), .Z(\_CLINT_io_rdata [11] ) );
BUF_X1 \CLINT/_1520_ ( .A(\CLINT/mtime [44] ), .Z(\CLINT/_0211_ ) );
BUF_X1 \CLINT/_1521_ ( .A(\CLINT/mtime [12] ), .Z(\CLINT/_0176_ ) );
BUF_X1 \CLINT/_1522_ ( .A(\CLINT/_0139_ ), .Z(\_CLINT_io_rdata [12] ) );
BUF_X1 \CLINT/_1523_ ( .A(\CLINT/mtime [45] ), .Z(\CLINT/_0212_ ) );
BUF_X1 \CLINT/_1524_ ( .A(\CLINT/mtime [13] ), .Z(\CLINT/_0177_ ) );
BUF_X1 \CLINT/_1525_ ( .A(\CLINT/_0140_ ), .Z(\_CLINT_io_rdata [13] ) );
BUF_X1 \CLINT/_1526_ ( .A(\CLINT/mtime [46] ), .Z(\CLINT/_0213_ ) );
BUF_X1 \CLINT/_1527_ ( .A(\CLINT/mtime [14] ), .Z(\CLINT/_0178_ ) );
BUF_X1 \CLINT/_1528_ ( .A(\CLINT/_0141_ ), .Z(\_CLINT_io_rdata [14] ) );
BUF_X1 \CLINT/_1529_ ( .A(\CLINT/mtime [47] ), .Z(\CLINT/_0214_ ) );
BUF_X1 \CLINT/_1530_ ( .A(\CLINT/mtime [15] ), .Z(\CLINT/_0179_ ) );
BUF_X1 \CLINT/_1531_ ( .A(\CLINT/_0142_ ), .Z(\_CLINT_io_rdata [15] ) );
BUF_X1 \CLINT/_1532_ ( .A(\CLINT/mtime [48] ), .Z(\CLINT/_0215_ ) );
BUF_X1 \CLINT/_1533_ ( .A(\CLINT/mtime [16] ), .Z(\CLINT/_0180_ ) );
BUF_X1 \CLINT/_1534_ ( .A(\CLINT/_0143_ ), .Z(\_CLINT_io_rdata [16] ) );
BUF_X1 \CLINT/_1535_ ( .A(\CLINT/mtime [49] ), .Z(\CLINT/_0216_ ) );
BUF_X1 \CLINT/_1536_ ( .A(\CLINT/mtime [17] ), .Z(\CLINT/_0181_ ) );
BUF_X1 \CLINT/_1537_ ( .A(\CLINT/_0144_ ), .Z(\_CLINT_io_rdata [17] ) );
BUF_X1 \CLINT/_1538_ ( .A(\CLINT/mtime [50] ), .Z(\CLINT/_0218_ ) );
BUF_X1 \CLINT/_1539_ ( .A(\CLINT/mtime [18] ), .Z(\CLINT/_0182_ ) );
BUF_X1 \CLINT/_1540_ ( .A(\CLINT/_0145_ ), .Z(\_CLINT_io_rdata [18] ) );
BUF_X1 \CLINT/_1541_ ( .A(\CLINT/mtime [51] ), .Z(\CLINT/_0219_ ) );
BUF_X1 \CLINT/_1542_ ( .A(\CLINT/mtime [19] ), .Z(\CLINT/_0183_ ) );
BUF_X1 \CLINT/_1543_ ( .A(\CLINT/_0146_ ), .Z(\_CLINT_io_rdata [19] ) );
BUF_X1 \CLINT/_1544_ ( .A(\CLINT/mtime [52] ), .Z(\CLINT/_0220_ ) );
BUF_X1 \CLINT/_1545_ ( .A(\CLINT/mtime [20] ), .Z(\CLINT/_0185_ ) );
BUF_X1 \CLINT/_1546_ ( .A(\CLINT/_0148_ ), .Z(\_CLINT_io_rdata [20] ) );
BUF_X1 \CLINT/_1547_ ( .A(\CLINT/mtime [53] ), .Z(\CLINT/_0221_ ) );
BUF_X1 \CLINT/_1548_ ( .A(\CLINT/mtime [21] ), .Z(\CLINT/_0186_ ) );
BUF_X1 \CLINT/_1549_ ( .A(\CLINT/_0149_ ), .Z(\_CLINT_io_rdata [21] ) );
BUF_X1 \CLINT/_1550_ ( .A(\CLINT/mtime [54] ), .Z(\CLINT/_0222_ ) );
BUF_X1 \CLINT/_1551_ ( .A(\CLINT/mtime [22] ), .Z(\CLINT/_0187_ ) );
BUF_X1 \CLINT/_1552_ ( .A(\CLINT/_0150_ ), .Z(\_CLINT_io_rdata [22] ) );
BUF_X1 \CLINT/_1553_ ( .A(\CLINT/mtime [55] ), .Z(\CLINT/_0223_ ) );
BUF_X1 \CLINT/_1554_ ( .A(\CLINT/mtime [23] ), .Z(\CLINT/_0188_ ) );
BUF_X1 \CLINT/_1555_ ( .A(\CLINT/_0151_ ), .Z(\_CLINT_io_rdata [23] ) );
BUF_X1 \CLINT/_1556_ ( .A(\CLINT/mtime [56] ), .Z(\CLINT/_0224_ ) );
BUF_X1 \CLINT/_1557_ ( .A(\CLINT/mtime [24] ), .Z(\CLINT/_0189_ ) );
BUF_X1 \CLINT/_1558_ ( .A(\CLINT/_0152_ ), .Z(\_CLINT_io_rdata [24] ) );
BUF_X1 \CLINT/_1559_ ( .A(\CLINT/mtime [57] ), .Z(\CLINT/_0225_ ) );
BUF_X1 \CLINT/_1560_ ( .A(\CLINT/mtime [25] ), .Z(\CLINT/_0190_ ) );
BUF_X1 \CLINT/_1561_ ( .A(\CLINT/_0153_ ), .Z(\_CLINT_io_rdata [25] ) );
BUF_X1 \CLINT/_1562_ ( .A(\CLINT/mtime [58] ), .Z(\CLINT/_0226_ ) );
BUF_X1 \CLINT/_1563_ ( .A(\CLINT/mtime [26] ), .Z(\CLINT/_0191_ ) );
BUF_X1 \CLINT/_1564_ ( .A(\CLINT/_0154_ ), .Z(\_CLINT_io_rdata [26] ) );
BUF_X1 \CLINT/_1565_ ( .A(\CLINT/mtime [59] ), .Z(\CLINT/_0227_ ) );
BUF_X1 \CLINT/_1566_ ( .A(\CLINT/mtime [27] ), .Z(\CLINT/_0192_ ) );
BUF_X1 \CLINT/_1567_ ( .A(\CLINT/_0155_ ), .Z(\_CLINT_io_rdata [27] ) );
BUF_X1 \CLINT/_1568_ ( .A(\CLINT/mtime [60] ), .Z(\CLINT/_0229_ ) );
BUF_X1 \CLINT/_1569_ ( .A(\CLINT/mtime [28] ), .Z(\CLINT/_0193_ ) );
BUF_X1 \CLINT/_1570_ ( .A(\CLINT/_0156_ ), .Z(\_CLINT_io_rdata [28] ) );
BUF_X1 \CLINT/_1571_ ( .A(\CLINT/mtime [61] ), .Z(\CLINT/_0230_ ) );
BUF_X1 \CLINT/_1572_ ( .A(\CLINT/mtime [29] ), .Z(\CLINT/_0194_ ) );
BUF_X1 \CLINT/_1573_ ( .A(\CLINT/_0157_ ), .Z(\_CLINT_io_rdata [29] ) );
BUF_X1 \CLINT/_1574_ ( .A(\CLINT/mtime [62] ), .Z(\CLINT/_0231_ ) );
BUF_X1 \CLINT/_1575_ ( .A(\CLINT/mtime [30] ), .Z(\CLINT/_0196_ ) );
BUF_X1 \CLINT/_1576_ ( .A(\CLINT/_0159_ ), .Z(\_CLINT_io_rdata [30] ) );
BUF_X1 \CLINT/_1577_ ( .A(\CLINT/mtime [63] ), .Z(\CLINT/_0232_ ) );
BUF_X1 \CLINT/_1578_ ( .A(\CLINT/mtime [31] ), .Z(\CLINT/_0197_ ) );
BUF_X1 \CLINT/_1579_ ( .A(\CLINT/_0160_ ), .Z(\_CLINT_io_rdata [31] ) );
BUF_X1 \CLINT/_1580_ ( .A(_AXI4Interconnect_io_fanOut_0_arvalid ), .Z(\CLINT/_0131_ ) );
BUF_X1 \CLINT/_1581_ ( .A(_AXI4Interconnect_io_fanOut_0_bready ), .Z(\CLINT/_0134_ ) );
BUF_X1 \CLINT/_1582_ ( .A(_AXI4Interconnect_io_fanOut_0_wvalid ), .Z(\CLINT/_0172_ ) );
BUF_X1 \CLINT/_1583_ ( .A(\CLINT/_0130_ ), .Z(_CLINT_io_arready ) );
BUF_X1 \CLINT/_1584_ ( .A(_AXI4Interconnect_io_fanOut_0_awvalid ), .Z(\CLINT/_0133_ ) );
BUF_X1 \CLINT/_1585_ ( .A(_AXI4Interconnect_io_fanOut_0_rready ), .Z(\CLINT/_0168_ ) );
BUF_X1 \CLINT/_1586_ ( .A(\CLINT/_0132_ ), .Z(_CLINT_io_awready ) );
BUF_X1 \CLINT/_1587_ ( .A(\CLINT/_0171_ ), .Z(_CLINT_io_wready ) );
BUF_X1 \CLINT/_1588_ ( .A(\CLINT/_0169_ ), .Z(\_CLINT_io_rresp [1] ) );
BUF_X1 \CLINT/_1589_ ( .A(\_AXI4Interconnect_io_fanOut_0_araddr [2] ), .Z(\CLINT/_0120_ ) );
BUF_X1 \CLINT/_1590_ ( .A(\CLINT/_0005_ ), .Z(\CLINT/_0743_ ) );
BUF_X1 \CLINT/_1591_ ( .A(\_AXI4Interconnect_io_fanOut_0_araddr [3] ), .Z(\CLINT/_0123_ ) );
BUF_X1 \CLINT/_1592_ ( .A(\CLINT/_0006_ ), .Z(\CLINT/_0744_ ) );
BUF_X1 \CLINT/_1593_ ( .A(\_AXI4Interconnect_io_fanOut_0_araddr [4] ), .Z(\CLINT/_0124_ ) );
BUF_X1 \CLINT/_1594_ ( .A(\CLINT/_0007_ ), .Z(\CLINT/_0745_ ) );
BUF_X1 \CLINT/_1595_ ( .A(\_AXI4Interconnect_io_fanOut_0_araddr [5] ), .Z(\CLINT/_0125_ ) );
BUF_X1 \CLINT/_1596_ ( .A(\CLINT/_0008_ ), .Z(\CLINT/_0746_ ) );
BUF_X1 \CLINT/_1597_ ( .A(\_AXI4Interconnect_io_fanOut_0_araddr [6] ), .Z(\CLINT/_0126_ ) );
BUF_X1 \CLINT/_1598_ ( .A(\CLINT/_0009_ ), .Z(\CLINT/_0747_ ) );
BUF_X1 \CLINT/_1599_ ( .A(\_AXI4Interconnect_io_fanOut_0_araddr [7] ), .Z(\CLINT/_0127_ ) );
BUF_X1 \CLINT/_1600_ ( .A(\CLINT/_0010_ ), .Z(\CLINT/_0748_ ) );
BUF_X1 \CLINT/_1601_ ( .A(\_AXI4Interconnect_io_fanOut_0_araddr [8] ), .Z(\CLINT/_0128_ ) );
BUF_X1 \CLINT/_1602_ ( .A(\CLINT/_0011_ ), .Z(\CLINT/_0749_ ) );
BUF_X1 \CLINT/_1603_ ( .A(\_AXI4Interconnect_io_fanOut_0_araddr [9] ), .Z(\CLINT/_0129_ ) );
BUF_X1 \CLINT/_1604_ ( .A(\CLINT/_0012_ ), .Z(\CLINT/_0750_ ) );
BUF_X1 \CLINT/_1605_ ( .A(\_AXI4Interconnect_io_fanOut_0_araddr [10] ), .Z(\CLINT/_0100_ ) );
BUF_X1 \CLINT/_1606_ ( .A(\CLINT/_0013_ ), .Z(\CLINT/_0751_ ) );
BUF_X1 \CLINT/_1607_ ( .A(\_AXI4Interconnect_io_fanOut_0_araddr [11] ), .Z(\CLINT/_0101_ ) );
BUF_X1 \CLINT/_1608_ ( .A(\CLINT/_0014_ ), .Z(\CLINT/_0752_ ) );
BUF_X1 \CLINT/_1609_ ( .A(\_AXI4Interconnect_io_fanOut_0_araddr [12] ), .Z(\CLINT/_0102_ ) );
BUF_X1 \CLINT/_1610_ ( .A(\CLINT/_0015_ ), .Z(\CLINT/_0753_ ) );
BUF_X1 \CLINT/_1611_ ( .A(\_AXI4Interconnect_io_fanOut_0_araddr [13] ), .Z(\CLINT/_0103_ ) );
BUF_X1 \CLINT/_1612_ ( .A(\CLINT/_0016_ ), .Z(\CLINT/_0754_ ) );
BUF_X1 \CLINT/_1613_ ( .A(\_AXI4Interconnect_io_fanOut_0_araddr [14] ), .Z(\CLINT/_0104_ ) );
BUF_X1 \CLINT/_1614_ ( .A(\CLINT/_0017_ ), .Z(\CLINT/_0755_ ) );
BUF_X1 \CLINT/_1615_ ( .A(\_AXI4Interconnect_io_fanOut_0_araddr [15] ), .Z(\CLINT/_0105_ ) );
BUF_X1 \CLINT/_1616_ ( .A(\CLINT/_0018_ ), .Z(\CLINT/_0756_ ) );
BUF_X1 \CLINT/_1617_ ( .A(\_AXI4Interconnect_io_fanOut_0_araddr [16] ), .Z(\CLINT/_0106_ ) );
BUF_X1 \CLINT/_1618_ ( .A(\CLINT/_0019_ ), .Z(\CLINT/_0757_ ) );
BUF_X1 \CLINT/_1619_ ( .A(\_AXI4Interconnect_io_fanOut_0_araddr [17] ), .Z(\CLINT/_0107_ ) );
BUF_X1 \CLINT/_1620_ ( .A(\CLINT/_0020_ ), .Z(\CLINT/_0758_ ) );
BUF_X1 \CLINT/_1621_ ( .A(\_AXI4Interconnect_io_fanOut_0_araddr [18] ), .Z(\CLINT/_0108_ ) );
BUF_X1 \CLINT/_1622_ ( .A(\CLINT/_0021_ ), .Z(\CLINT/_0759_ ) );
BUF_X1 \CLINT/_1623_ ( .A(\_AXI4Interconnect_io_fanOut_0_araddr [19] ), .Z(\CLINT/_0109_ ) );
BUF_X1 \CLINT/_1624_ ( .A(\CLINT/_0022_ ), .Z(\CLINT/_0760_ ) );
BUF_X1 \CLINT/_1625_ ( .A(\_AXI4Interconnect_io_fanOut_0_araddr [20] ), .Z(\CLINT/_0110_ ) );
BUF_X1 \CLINT/_1626_ ( .A(\CLINT/_0023_ ), .Z(\CLINT/_0761_ ) );
BUF_X1 \CLINT/_1627_ ( .A(\_AXI4Interconnect_io_fanOut_0_araddr [21] ), .Z(\CLINT/_0111_ ) );
BUF_X1 \CLINT/_1628_ ( .A(\CLINT/_0024_ ), .Z(\CLINT/_0762_ ) );
BUF_X1 \CLINT/_1629_ ( .A(\_AXI4Interconnect_io_fanOut_0_araddr [22] ), .Z(\CLINT/_0112_ ) );
BUF_X1 \CLINT/_1630_ ( .A(\CLINT/_0025_ ), .Z(\CLINT/_0763_ ) );
BUF_X1 \CLINT/_1631_ ( .A(\_AXI4Interconnect_io_fanOut_0_araddr [23] ), .Z(\CLINT/_0113_ ) );
BUF_X1 \CLINT/_1632_ ( .A(\CLINT/_0026_ ), .Z(\CLINT/_0764_ ) );
BUF_X1 \CLINT/_1633_ ( .A(\_AXI4Interconnect_io_fanOut_0_araddr [24] ), .Z(\CLINT/_0114_ ) );
BUF_X1 \CLINT/_1634_ ( .A(\CLINT/_0027_ ), .Z(\CLINT/_0765_ ) );
BUF_X1 \CLINT/_1635_ ( .A(\_AXI4Interconnect_io_fanOut_0_araddr [25] ), .Z(\CLINT/_0115_ ) );
BUF_X1 \CLINT/_1636_ ( .A(\CLINT/_0028_ ), .Z(\CLINT/_0766_ ) );
BUF_X1 \CLINT/_1637_ ( .A(\_AXI4Interconnect_io_fanOut_0_araddr [26] ), .Z(\CLINT/_0116_ ) );
BUF_X1 \CLINT/_1638_ ( .A(\CLINT/_0029_ ), .Z(\CLINT/_0767_ ) );
BUF_X1 \CLINT/_1639_ ( .A(\_AXI4Interconnect_io_fanOut_0_araddr [27] ), .Z(\CLINT/_0117_ ) );
BUF_X1 \CLINT/_1640_ ( .A(\CLINT/_0030_ ), .Z(\CLINT/_0768_ ) );
BUF_X1 \CLINT/_1641_ ( .A(\_AXI4Interconnect_io_fanOut_0_araddr [28] ), .Z(\CLINT/_0118_ ) );
BUF_X1 \CLINT/_1642_ ( .A(\CLINT/_0031_ ), .Z(\CLINT/_0769_ ) );
BUF_X1 \CLINT/_1643_ ( .A(\_AXI4Interconnect_io_fanOut_0_araddr [29] ), .Z(\CLINT/_0119_ ) );
BUF_X1 \CLINT/_1644_ ( .A(\CLINT/_0032_ ), .Z(\CLINT/_0770_ ) );
BUF_X1 \CLINT/_1645_ ( .A(\_AXI4Interconnect_io_fanOut_0_araddr [30] ), .Z(\CLINT/_0121_ ) );
BUF_X1 \CLINT/_1646_ ( .A(\CLINT/_0033_ ), .Z(\CLINT/_0771_ ) );
BUF_X1 \CLINT/_1647_ ( .A(\_AXI4Interconnect_io_fanOut_0_araddr [31] ), .Z(\CLINT/_0122_ ) );
BUF_X1 \CLINT/_1648_ ( .A(\CLINT/_0034_ ), .Z(\CLINT/_0772_ ) );
BUF_X1 \CLINT/_1649_ ( .A(\CLINT/_0003_ ), .Z(\CLINT/_0741_ ) );
BUF_X1 \CLINT/_1650_ ( .A(\CLINT/_0004_ ), .Z(\CLINT/_0742_ ) );
BUF_X1 \CLINT/_1651_ ( .A(\CLINT/_0035_ ), .Z(\CLINT/_0773_ ) );
BUF_X1 \CLINT/_1652_ ( .A(\CLINT/_0581_ ), .Z(\CLINT/_0002_ ) );
BUF_X1 \CLINT/_1653_ ( .A(\CLINT/_0036_ ), .Z(\CLINT/_0774_ ) );
BUF_X1 \CLINT/_1654_ ( .A(\CLINT/_0037_ ), .Z(\CLINT/_0775_ ) );
BUF_X1 \CLINT/_1655_ ( .A(\CLINT/_0038_ ), .Z(\CLINT/_0776_ ) );
BUF_X1 \CLINT/_1656_ ( .A(\CLINT/_0039_ ), .Z(\CLINT/_0777_ ) );
BUF_X1 \CLINT/_1657_ ( .A(\CLINT/_0040_ ), .Z(\CLINT/_0778_ ) );
BUF_X1 \CLINT/_1658_ ( .A(\CLINT/_0041_ ), .Z(\CLINT/_0779_ ) );
BUF_X1 \CLINT/_1659_ ( .A(\CLINT/_0042_ ), .Z(\CLINT/_0780_ ) );
BUF_X1 \CLINT/_1660_ ( .A(\CLINT/_0043_ ), .Z(\CLINT/_0781_ ) );
BUF_X1 \CLINT/_1661_ ( .A(\CLINT/_0044_ ), .Z(\CLINT/_0782_ ) );
BUF_X1 \CLINT/_1662_ ( .A(\CLINT/_0045_ ), .Z(\CLINT/_0783_ ) );
BUF_X1 \CLINT/_1663_ ( .A(\CLINT/_0046_ ), .Z(\CLINT/_0784_ ) );
BUF_X1 \CLINT/_1664_ ( .A(\CLINT/_0047_ ), .Z(\CLINT/_0785_ ) );
BUF_X1 \CLINT/_1665_ ( .A(\CLINT/_0048_ ), .Z(\CLINT/_0786_ ) );
BUF_X1 \CLINT/_1666_ ( .A(\CLINT/_0049_ ), .Z(\CLINT/_0787_ ) );
BUF_X1 \CLINT/_1667_ ( .A(\CLINT/_0050_ ), .Z(\CLINT/_0788_ ) );
BUF_X1 \CLINT/_1668_ ( .A(\CLINT/_0051_ ), .Z(\CLINT/_0789_ ) );
BUF_X1 \CLINT/_1669_ ( .A(\CLINT/_0052_ ), .Z(\CLINT/_0790_ ) );
BUF_X1 \CLINT/_1670_ ( .A(\CLINT/_0053_ ), .Z(\CLINT/_0791_ ) );
BUF_X1 \CLINT/_1671_ ( .A(\CLINT/_0054_ ), .Z(\CLINT/_0792_ ) );
BUF_X1 \CLINT/_1672_ ( .A(\CLINT/_0055_ ), .Z(\CLINT/_0793_ ) );
BUF_X1 \CLINT/_1673_ ( .A(\CLINT/_0056_ ), .Z(\CLINT/_0794_ ) );
BUF_X1 \CLINT/_1674_ ( .A(\CLINT/_0057_ ), .Z(\CLINT/_0795_ ) );
BUF_X1 \CLINT/_1675_ ( .A(\CLINT/_0058_ ), .Z(\CLINT/_0796_ ) );
BUF_X1 \CLINT/_1676_ ( .A(\CLINT/_0059_ ), .Z(\CLINT/_0797_ ) );
BUF_X1 \CLINT/_1677_ ( .A(\CLINT/_0060_ ), .Z(\CLINT/_0798_ ) );
BUF_X1 \CLINT/_1678_ ( .A(\CLINT/_0061_ ), .Z(\CLINT/_0799_ ) );
BUF_X1 \CLINT/_1679_ ( .A(\CLINT/_0062_ ), .Z(\CLINT/_0800_ ) );
BUF_X1 \CLINT/_1680_ ( .A(\CLINT/_0063_ ), .Z(\CLINT/_0801_ ) );
BUF_X1 \CLINT/_1681_ ( .A(\CLINT/_0064_ ), .Z(\CLINT/_0802_ ) );
BUF_X1 \CLINT/_1682_ ( .A(\CLINT/_0065_ ), .Z(\CLINT/_0803_ ) );
BUF_X1 \CLINT/_1683_ ( .A(\CLINT/_0066_ ), .Z(\CLINT/_0804_ ) );
BUF_X1 \CLINT/_1684_ ( .A(\CLINT/_0067_ ), .Z(\CLINT/_0805_ ) );
BUF_X1 \CLINT/_1685_ ( .A(\CLINT/_0068_ ), .Z(\CLINT/_0806_ ) );
BUF_X1 \CLINT/_1686_ ( .A(\CLINT/_0069_ ), .Z(\CLINT/_0807_ ) );
BUF_X1 \CLINT/_1687_ ( .A(\CLINT/_0070_ ), .Z(\CLINT/_0808_ ) );
BUF_X1 \CLINT/_1688_ ( .A(\CLINT/_0071_ ), .Z(\CLINT/_0809_ ) );
BUF_X1 \CLINT/_1689_ ( .A(\CLINT/_0072_ ), .Z(\CLINT/_0810_ ) );
BUF_X1 \CLINT/_1690_ ( .A(\CLINT/_0073_ ), .Z(\CLINT/_0811_ ) );
BUF_X1 \CLINT/_1691_ ( .A(\CLINT/_0074_ ), .Z(\CLINT/_0812_ ) );
BUF_X1 \CLINT/_1692_ ( .A(\CLINT/_0075_ ), .Z(\CLINT/_0813_ ) );
BUF_X1 \CLINT/_1693_ ( .A(\CLINT/_0076_ ), .Z(\CLINT/_0814_ ) );
BUF_X1 \CLINT/_1694_ ( .A(\CLINT/_0077_ ), .Z(\CLINT/_0815_ ) );
BUF_X1 \CLINT/_1695_ ( .A(\CLINT/_0078_ ), .Z(\CLINT/_0816_ ) );
BUF_X1 \CLINT/_1696_ ( .A(\CLINT/_0079_ ), .Z(\CLINT/_0817_ ) );
BUF_X1 \CLINT/_1697_ ( .A(\CLINT/_0080_ ), .Z(\CLINT/_0818_ ) );
BUF_X1 \CLINT/_1698_ ( .A(\CLINT/_0081_ ), .Z(\CLINT/_0819_ ) );
BUF_X1 \CLINT/_1699_ ( .A(\CLINT/_0082_ ), .Z(\CLINT/_0820_ ) );
BUF_X1 \CLINT/_1700_ ( .A(\CLINT/_0083_ ), .Z(\CLINT/_0821_ ) );
BUF_X1 \CLINT/_1701_ ( .A(\CLINT/_0084_ ), .Z(\CLINT/_0822_ ) );
BUF_X1 \CLINT/_1702_ ( .A(\CLINT/_0085_ ), .Z(\CLINT/_0823_ ) );
BUF_X1 \CLINT/_1703_ ( .A(\CLINT/_0086_ ), .Z(\CLINT/_0824_ ) );
BUF_X1 \CLINT/_1704_ ( .A(\CLINT/_0087_ ), .Z(\CLINT/_0825_ ) );
BUF_X1 \CLINT/_1705_ ( .A(\CLINT/_0088_ ), .Z(\CLINT/_0826_ ) );
BUF_X1 \CLINT/_1706_ ( .A(\CLINT/_0089_ ), .Z(\CLINT/_0827_ ) );
BUF_X1 \CLINT/_1707_ ( .A(\CLINT/_0090_ ), .Z(\CLINT/_0828_ ) );
BUF_X1 \CLINT/_1708_ ( .A(\CLINT/_0091_ ), .Z(\CLINT/_0829_ ) );
BUF_X1 \CLINT/_1709_ ( .A(\CLINT/_0092_ ), .Z(\CLINT/_0830_ ) );
BUF_X1 \CLINT/_1710_ ( .A(\CLINT/_0093_ ), .Z(\CLINT/_0831_ ) );
BUF_X1 \CLINT/_1711_ ( .A(\CLINT/_0094_ ), .Z(\CLINT/_0832_ ) );
BUF_X1 \CLINT/_1712_ ( .A(\CLINT/_0095_ ), .Z(\CLINT/_0833_ ) );
BUF_X1 \CLINT/_1713_ ( .A(\CLINT/_0096_ ), .Z(\CLINT/_0834_ ) );
BUF_X1 \CLINT/_1714_ ( .A(\CLINT/_0097_ ), .Z(\CLINT/_0835_ ) );
BUF_X1 \CLINT/_1715_ ( .A(\CLINT/_0098_ ), .Z(\CLINT/_0836_ ) );
BUF_X1 \CLINT/_1716_ ( .A(\CLINT/_0099_ ), .Z(\CLINT/_0837_ ) );
AND2_X1 \EXU/_1643_ ( .A1(\EXU/_1215_ ), .A2(\EXU/_1216_ ), .ZN(\EXU/_0842_ ) );
INV_X1 \EXU/_1644_ ( .A(\EXU/_1215_ ), .ZN(\EXU/_1101_ ) );
AND2_X1 \EXU/_1645_ ( .A1(\EXU/_1101_ ), .A2(\EXU/_1216_ ), .ZN(\EXU/_0594_ ) );
NOR2_X1 \EXU/_1646_ ( .A1(\EXU/_1101_ ), .A2(\EXU/_1216_ ), .ZN(\EXU/_0561_ ) );
NOR2_X1 \EXU/_1647_ ( .A1(\EXU/_1215_ ), .A2(\EXU/_1216_ ), .ZN(\EXU/_0775_ ) );
MUX2_X1 \EXU/_1648_ ( .A(\EXU/_0459_ ), .B(\EXU/_0427_ ), .S(fanout_net_10 ), .Z(\EXU/_0069_ ) );
MUX2_X1 \EXU/_1649_ ( .A(\EXU/_0470_ ), .B(\EXU/_0438_ ), .S(fanout_net_10 ), .Z(\EXU/_0080_ ) );
MUX2_X1 \EXU/_1650_ ( .A(\EXU/_0481_ ), .B(\EXU/_0449_ ), .S(fanout_net_10 ), .Z(\EXU/_0091_ ) );
MUX2_X1 \EXU/_1651_ ( .A(\EXU/_0484_ ), .B(\EXU/_0452_ ), .S(fanout_net_10 ), .Z(\EXU/_0094_ ) );
MUX2_X1 \EXU/_1652_ ( .A(\EXU/_0485_ ), .B(\EXU/_0453_ ), .S(fanout_net_10 ), .Z(\EXU/_0095_ ) );
MUX2_X1 \EXU/_1653_ ( .A(\EXU/_0486_ ), .B(\EXU/_0454_ ), .S(fanout_net_10 ), .Z(\EXU/_0096_ ) );
MUX2_X1 \EXU/_1654_ ( .A(\EXU/_0487_ ), .B(\EXU/_0455_ ), .S(fanout_net_10 ), .Z(\EXU/_0097_ ) );
MUX2_X1 \EXU/_1655_ ( .A(\EXU/_0488_ ), .B(\EXU/_0456_ ), .S(fanout_net_10 ), .Z(\EXU/_0098_ ) );
MUX2_X1 \EXU/_1656_ ( .A(\EXU/_0489_ ), .B(\EXU/_0457_ ), .S(fanout_net_10 ), .Z(\EXU/_0099_ ) );
MUX2_X1 \EXU/_1657_ ( .A(\EXU/_0490_ ), .B(\EXU/_0458_ ), .S(fanout_net_10 ), .Z(\EXU/_0100_ ) );
MUX2_X1 \EXU/_1658_ ( .A(\EXU/_0460_ ), .B(\EXU/_0428_ ), .S(fanout_net_10 ), .Z(\EXU/_0070_ ) );
MUX2_X1 \EXU/_1659_ ( .A(\EXU/_0461_ ), .B(\EXU/_0429_ ), .S(fanout_net_10 ), .Z(\EXU/_0071_ ) );
MUX2_X1 \EXU/_1660_ ( .A(\EXU/_0462_ ), .B(\EXU/_0430_ ), .S(fanout_net_10 ), .Z(\EXU/_0072_ ) );
MUX2_X1 \EXU/_1661_ ( .A(\EXU/_0463_ ), .B(\EXU/_0431_ ), .S(fanout_net_10 ), .Z(\EXU/_0073_ ) );
MUX2_X1 \EXU/_1662_ ( .A(\EXU/_0464_ ), .B(\EXU/_0432_ ), .S(fanout_net_10 ), .Z(\EXU/_0074_ ) );
MUX2_X1 \EXU/_1663_ ( .A(\EXU/_0465_ ), .B(\EXU/_0433_ ), .S(fanout_net_10 ), .Z(\EXU/_0075_ ) );
MUX2_X1 \EXU/_1664_ ( .A(\EXU/_0466_ ), .B(\EXU/_0434_ ), .S(fanout_net_10 ), .Z(\EXU/_0076_ ) );
MUX2_X1 \EXU/_1665_ ( .A(\EXU/_0467_ ), .B(\EXU/_0435_ ), .S(fanout_net_10 ), .Z(\EXU/_0077_ ) );
MUX2_X1 \EXU/_1666_ ( .A(\EXU/_0468_ ), .B(\EXU/_0436_ ), .S(fanout_net_10 ), .Z(\EXU/_0078_ ) );
MUX2_X1 \EXU/_1667_ ( .A(\EXU/_0469_ ), .B(\EXU/_0437_ ), .S(fanout_net_10 ), .Z(\EXU/_0079_ ) );
MUX2_X1 \EXU/_1668_ ( .A(\EXU/_0471_ ), .B(\EXU/_0439_ ), .S(fanout_net_10 ), .Z(\EXU/_0081_ ) );
MUX2_X1 \EXU/_1669_ ( .A(\EXU/_0472_ ), .B(\EXU/_0440_ ), .S(fanout_net_10 ), .Z(\EXU/_0082_ ) );
MUX2_X1 \EXU/_1670_ ( .A(\EXU/_0473_ ), .B(\EXU/_0441_ ), .S(fanout_net_10 ), .Z(\EXU/_0083_ ) );
MUX2_X1 \EXU/_1671_ ( .A(\EXU/_0474_ ), .B(\EXU/_0442_ ), .S(fanout_net_10 ), .Z(\EXU/_0084_ ) );
MUX2_X1 \EXU/_1672_ ( .A(\EXU/_0475_ ), .B(\EXU/_0443_ ), .S(fanout_net_10 ), .Z(\EXU/_0085_ ) );
MUX2_X1 \EXU/_1673_ ( .A(\EXU/_0476_ ), .B(\EXU/_0444_ ), .S(fanout_net_10 ), .Z(\EXU/_0086_ ) );
MUX2_X1 \EXU/_1674_ ( .A(\EXU/_0477_ ), .B(\EXU/_0445_ ), .S(fanout_net_10 ), .Z(\EXU/_0087_ ) );
MUX2_X1 \EXU/_1675_ ( .A(\EXU/_0478_ ), .B(\EXU/_0446_ ), .S(fanout_net_10 ), .Z(\EXU/_0088_ ) );
MUX2_X1 \EXU/_1676_ ( .A(\EXU/_0479_ ), .B(\EXU/_0447_ ), .S(fanout_net_10 ), .Z(\EXU/_0089_ ) );
MUX2_X1 \EXU/_1677_ ( .A(\EXU/_0480_ ), .B(\EXU/_0448_ ), .S(fanout_net_10 ), .Z(\EXU/_0090_ ) );
MUX2_X1 \EXU/_1678_ ( .A(\EXU/_0482_ ), .B(\EXU/_0450_ ), .S(\EXU/_0381_ ), .Z(\EXU/_0092_ ) );
MUX2_X1 \EXU/_1679_ ( .A(\EXU/_0483_ ), .B(\EXU/_0451_ ), .S(\EXU/_0381_ ), .Z(\EXU/_0093_ ) );
AND3_X1 \EXU/_1680_ ( .A1(\EXU/_1215_ ), .A2(\EXU/_1216_ ), .A3(\EXU/_0391_ ), .ZN(\EXU/_0101_ ) );
AND3_X1 \EXU/_1681_ ( .A1(\EXU/_1215_ ), .A2(\EXU/_1216_ ), .A3(\EXU/_0392_ ), .ZN(\EXU/_0102_ ) );
AND3_X1 \EXU/_1682_ ( .A1(\EXU/_1215_ ), .A2(\EXU/_1216_ ), .A3(\EXU/_0393_ ), .ZN(\EXU/_0103_ ) );
MUX2_X1 \EXU/_1683_ ( .A(\EXU/_0459_ ), .B(\EXU/_0491_ ), .S(fanout_net_11 ), .Z(\EXU/_0104_ ) );
MUX2_X1 \EXU/_1684_ ( .A(\EXU/_0470_ ), .B(\EXU/_0502_ ), .S(fanout_net_11 ), .Z(\EXU/_0115_ ) );
MUX2_X1 \EXU/_1685_ ( .A(\EXU/_0481_ ), .B(\EXU/_0513_ ), .S(fanout_net_11 ), .Z(\EXU/_0126_ ) );
MUX2_X1 \EXU/_1686_ ( .A(\EXU/_0484_ ), .B(\EXU/_0516_ ), .S(fanout_net_11 ), .Z(\EXU/_0129_ ) );
MUX2_X1 \EXU/_1687_ ( .A(\EXU/_0485_ ), .B(\EXU/_0517_ ), .S(fanout_net_11 ), .Z(\EXU/_0130_ ) );
MUX2_X1 \EXU/_1688_ ( .A(\EXU/_0486_ ), .B(\EXU/_0518_ ), .S(fanout_net_11 ), .Z(\EXU/_0131_ ) );
MUX2_X1 \EXU/_1689_ ( .A(\EXU/_0487_ ), .B(\EXU/_0519_ ), .S(fanout_net_11 ), .Z(\EXU/_0132_ ) );
MUX2_X1 \EXU/_1690_ ( .A(\EXU/_0488_ ), .B(\EXU/_0520_ ), .S(fanout_net_11 ), .Z(\EXU/_0133_ ) );
MUX2_X1 \EXU/_1691_ ( .A(\EXU/_0489_ ), .B(\EXU/_0521_ ), .S(fanout_net_11 ), .Z(\EXU/_0134_ ) );
MUX2_X1 \EXU/_1692_ ( .A(\EXU/_0490_ ), .B(\EXU/_0522_ ), .S(fanout_net_11 ), .Z(\EXU/_0135_ ) );
MUX2_X1 \EXU/_1693_ ( .A(\EXU/_0460_ ), .B(\EXU/_0492_ ), .S(fanout_net_11 ), .Z(\EXU/_0105_ ) );
MUX2_X1 \EXU/_1694_ ( .A(\EXU/_0461_ ), .B(\EXU/_0493_ ), .S(fanout_net_11 ), .Z(\EXU/_0106_ ) );
MUX2_X1 \EXU/_1695_ ( .A(\EXU/_0462_ ), .B(\EXU/_0494_ ), .S(fanout_net_11 ), .Z(\EXU/_0107_ ) );
MUX2_X1 \EXU/_1696_ ( .A(\EXU/_0463_ ), .B(\EXU/_0495_ ), .S(fanout_net_11 ), .Z(\EXU/_0108_ ) );
MUX2_X1 \EXU/_1697_ ( .A(\EXU/_0464_ ), .B(\EXU/_0496_ ), .S(fanout_net_11 ), .Z(\EXU/_0109_ ) );
MUX2_X1 \EXU/_1698_ ( .A(\EXU/_0465_ ), .B(\EXU/_0497_ ), .S(fanout_net_11 ), .Z(\EXU/_0110_ ) );
MUX2_X1 \EXU/_1699_ ( .A(\EXU/_0466_ ), .B(\EXU/_0498_ ), .S(fanout_net_11 ), .Z(\EXU/_0111_ ) );
MUX2_X1 \EXU/_1700_ ( .A(\EXU/_0467_ ), .B(\EXU/_0499_ ), .S(fanout_net_11 ), .Z(\EXU/_0112_ ) );
MUX2_X1 \EXU/_1701_ ( .A(\EXU/_0468_ ), .B(\EXU/_0500_ ), .S(fanout_net_11 ), .Z(\EXU/_0113_ ) );
MUX2_X1 \EXU/_1702_ ( .A(\EXU/_0469_ ), .B(\EXU/_0501_ ), .S(fanout_net_11 ), .Z(\EXU/_0114_ ) );
MUX2_X1 \EXU/_1703_ ( .A(\EXU/_0471_ ), .B(\EXU/_0503_ ), .S(fanout_net_11 ), .Z(\EXU/_0116_ ) );
MUX2_X1 \EXU/_1704_ ( .A(\EXU/_0472_ ), .B(\EXU/_0504_ ), .S(fanout_net_11 ), .Z(\EXU/_0117_ ) );
MUX2_X1 \EXU/_1705_ ( .A(\EXU/_0473_ ), .B(\EXU/_0505_ ), .S(fanout_net_11 ), .Z(\EXU/_0118_ ) );
MUX2_X1 \EXU/_1706_ ( .A(\EXU/_0474_ ), .B(\EXU/_0506_ ), .S(fanout_net_11 ), .Z(\EXU/_0119_ ) );
MUX2_X1 \EXU/_1707_ ( .A(\EXU/_0475_ ), .B(\EXU/_0507_ ), .S(fanout_net_11 ), .Z(\EXU/_0120_ ) );
MUX2_X1 \EXU/_1708_ ( .A(\EXU/_0476_ ), .B(\EXU/_0508_ ), .S(fanout_net_11 ), .Z(\EXU/_0121_ ) );
MUX2_X1 \EXU/_1709_ ( .A(\EXU/_0477_ ), .B(\EXU/_0509_ ), .S(fanout_net_11 ), .Z(\EXU/_0122_ ) );
MUX2_X1 \EXU/_1710_ ( .A(\EXU/_0478_ ), .B(\EXU/_0510_ ), .S(fanout_net_11 ), .Z(\EXU/_0123_ ) );
MUX2_X1 \EXU/_1711_ ( .A(\EXU/_0479_ ), .B(\EXU/_0511_ ), .S(fanout_net_11 ), .Z(\EXU/_0124_ ) );
MUX2_X1 \EXU/_1712_ ( .A(\EXU/_0480_ ), .B(\EXU/_0512_ ), .S(fanout_net_11 ), .Z(\EXU/_0125_ ) );
MUX2_X1 \EXU/_1713_ ( .A(\EXU/_0482_ ), .B(\EXU/_0514_ ), .S(\EXU/_0394_ ), .Z(\EXU/_0127_ ) );
MUX2_X1 \EXU/_1714_ ( .A(\EXU/_0483_ ), .B(\EXU/_0515_ ), .S(\EXU/_0394_ ), .Z(\EXU/_0128_ ) );
INV_X1 \EXU/_1715_ ( .A(\EXU/_0382_ ), .ZN(\EXU/_1102_ ) );
NOR2_X1 \EXU/_1716_ ( .A1(\EXU/_1102_ ), .A2(\EXU/_0383_ ), .ZN(\EXU/_1103_ ) );
BUF_X4 \EXU/_1717_ ( .A(\EXU/_1103_ ), .Z(\EXU/_1104_ ) );
NAND2_X1 \EXU/_1718_ ( .A1(\EXU/_1104_ ), .A2(\EXU/_0395_ ), .ZN(\EXU/_1105_ ) );
NOR2_X1 \EXU/_1719_ ( .A1(\EXU/_0382_ ), .A2(\EXU/_0383_ ), .ZN(\EXU/_1106_ ) );
BUF_X4 \EXU/_1720_ ( .A(\EXU/_1106_ ), .Z(\EXU/_1107_ ) );
NAND2_X1 \EXU/_1721_ ( .A1(\EXU/_1107_ ), .A2(\EXU/_0527_ ), .ZN(\EXU/_1108_ ) );
NAND2_X1 \EXU/_1722_ ( .A1(\EXU/_1105_ ), .A2(\EXU/_1108_ ), .ZN(\EXU/_0349_ ) );
NAND2_X1 \EXU/_1723_ ( .A1(\EXU/_1104_ ), .A2(\EXU/_0406_ ), .ZN(\EXU/_1109_ ) );
NAND2_X1 \EXU/_1724_ ( .A1(\EXU/_1107_ ), .A2(\EXU/_0538_ ), .ZN(\EXU/_1110_ ) );
NAND2_X1 \EXU/_1725_ ( .A1(\EXU/_1109_ ), .A2(\EXU/_1110_ ), .ZN(\EXU/_0360_ ) );
NOR3_X1 \EXU/_1726_ ( .A1(\EXU/_0382_ ), .A2(\EXU/_0383_ ), .A3(\EXU/_0549_ ), .ZN(\EXU/_1111_ ) );
INV_X1 \EXU/_1727_ ( .A(\EXU/_0417_ ), .ZN(\EXU/_1112_ ) );
AOI21_X1 \EXU/_1728_ ( .A(\EXU/_1111_ ), .B1(\EXU/_1112_ ), .B2(\EXU/_1104_ ), .ZN(\EXU/_0371_ ) );
NAND2_X1 \EXU/_1729_ ( .A1(\EXU/_1104_ ), .A2(\EXU/_0420_ ), .ZN(\EXU/_1113_ ) );
NAND2_X1 \EXU/_1730_ ( .A1(\EXU/_1107_ ), .A2(\EXU/_0552_ ), .ZN(\EXU/_1114_ ) );
NAND2_X1 \EXU/_1731_ ( .A1(\EXU/_1113_ ), .A2(\EXU/_1114_ ), .ZN(\EXU/_0374_ ) );
NAND2_X1 \EXU/_1732_ ( .A1(\EXU/_1104_ ), .A2(\EXU/_0421_ ), .ZN(\EXU/_1115_ ) );
NAND2_X1 \EXU/_1733_ ( .A1(\EXU/_1107_ ), .A2(\EXU/_0553_ ), .ZN(\EXU/_1116_ ) );
NAND2_X1 \EXU/_1734_ ( .A1(\EXU/_1115_ ), .A2(\EXU/_1116_ ), .ZN(\EXU/_0375_ ) );
NAND2_X1 \EXU/_1735_ ( .A1(\EXU/_1104_ ), .A2(\EXU/_0422_ ), .ZN(\EXU/_1117_ ) );
NAND2_X1 \EXU/_1736_ ( .A1(\EXU/_1107_ ), .A2(\EXU/_0554_ ), .ZN(\EXU/_1118_ ) );
NAND2_X1 \EXU/_1737_ ( .A1(\EXU/_1117_ ), .A2(\EXU/_1118_ ), .ZN(\EXU/_0376_ ) );
NAND2_X1 \EXU/_1738_ ( .A1(\EXU/_1104_ ), .A2(\EXU/_0423_ ), .ZN(\EXU/_1119_ ) );
NAND2_X1 \EXU/_1739_ ( .A1(\EXU/_1107_ ), .A2(\EXU/_0555_ ), .ZN(\EXU/_1120_ ) );
NAND2_X1 \EXU/_1740_ ( .A1(\EXU/_1119_ ), .A2(\EXU/_1120_ ), .ZN(\EXU/_0377_ ) );
NAND2_X1 \EXU/_1741_ ( .A1(\EXU/_1104_ ), .A2(\EXU/_0424_ ), .ZN(\EXU/_1121_ ) );
NAND2_X1 \EXU/_1742_ ( .A1(\EXU/_1107_ ), .A2(\EXU/_0556_ ), .ZN(\EXU/_1122_ ) );
NAND2_X1 \EXU/_1743_ ( .A1(\EXU/_1121_ ), .A2(\EXU/_1122_ ), .ZN(\EXU/_0378_ ) );
NAND2_X1 \EXU/_1744_ ( .A1(\EXU/_1104_ ), .A2(\EXU/_0425_ ), .ZN(\EXU/_1123_ ) );
NAND2_X1 \EXU/_1745_ ( .A1(\EXU/_1107_ ), .A2(\EXU/_0557_ ), .ZN(\EXU/_1124_ ) );
NAND2_X1 \EXU/_1746_ ( .A1(\EXU/_1123_ ), .A2(\EXU/_1124_ ), .ZN(\EXU/_0379_ ) );
NAND2_X1 \EXU/_1747_ ( .A1(\EXU/_1104_ ), .A2(\EXU/_0426_ ), .ZN(\EXU/_1125_ ) );
NAND2_X1 \EXU/_1748_ ( .A1(\EXU/_1107_ ), .A2(\EXU/_0558_ ), .ZN(\EXU/_1126_ ) );
NAND2_X1 \EXU/_1749_ ( .A1(\EXU/_1125_ ), .A2(\EXU/_1126_ ), .ZN(\EXU/_0380_ ) );
BUF_X4 \EXU/_1750_ ( .A(\EXU/_1103_ ), .Z(\EXU/_1127_ ) );
NAND2_X1 \EXU/_1751_ ( .A1(\EXU/_1127_ ), .A2(\EXU/_0396_ ), .ZN(\EXU/_1128_ ) );
NAND2_X1 \EXU/_1752_ ( .A1(\EXU/_1107_ ), .A2(\EXU/_0528_ ), .ZN(\EXU/_1129_ ) );
NAND2_X1 \EXU/_1753_ ( .A1(\EXU/_1128_ ), .A2(\EXU/_1129_ ), .ZN(\EXU/_0350_ ) );
NAND2_X1 \EXU/_1754_ ( .A1(\EXU/_1127_ ), .A2(\EXU/_0397_ ), .ZN(\EXU/_1130_ ) );
BUF_X4 \EXU/_1755_ ( .A(\EXU/_1106_ ), .Z(\EXU/_1131_ ) );
NAND2_X1 \EXU/_1756_ ( .A1(\EXU/_1131_ ), .A2(\EXU/_0529_ ), .ZN(\EXU/_1132_ ) );
NAND2_X1 \EXU/_1757_ ( .A1(\EXU/_1130_ ), .A2(\EXU/_1132_ ), .ZN(\EXU/_0351_ ) );
NAND2_X1 \EXU/_1758_ ( .A1(\EXU/_1127_ ), .A2(\EXU/_0398_ ), .ZN(\EXU/_1133_ ) );
NAND2_X1 \EXU/_1759_ ( .A1(\EXU/_1131_ ), .A2(\EXU/_0530_ ), .ZN(\EXU/_1134_ ) );
NAND2_X1 \EXU/_1760_ ( .A1(\EXU/_1133_ ), .A2(\EXU/_1134_ ), .ZN(\EXU/_0352_ ) );
NAND2_X1 \EXU/_1761_ ( .A1(\EXU/_1127_ ), .A2(\EXU/_0399_ ), .ZN(\EXU/_1135_ ) );
NAND2_X1 \EXU/_1762_ ( .A1(\EXU/_1131_ ), .A2(\EXU/_0531_ ), .ZN(\EXU/_1136_ ) );
NAND2_X1 \EXU/_1763_ ( .A1(\EXU/_1135_ ), .A2(\EXU/_1136_ ), .ZN(\EXU/_0353_ ) );
NAND2_X1 \EXU/_1764_ ( .A1(\EXU/_1127_ ), .A2(\EXU/_0400_ ), .ZN(\EXU/_1137_ ) );
NAND2_X1 \EXU/_1765_ ( .A1(\EXU/_1131_ ), .A2(\EXU/_0532_ ), .ZN(\EXU/_1138_ ) );
NAND2_X1 \EXU/_1766_ ( .A1(\EXU/_1137_ ), .A2(\EXU/_1138_ ), .ZN(\EXU/_0354_ ) );
NAND2_X1 \EXU/_1767_ ( .A1(\EXU/_1127_ ), .A2(\EXU/_0401_ ), .ZN(\EXU/_1139_ ) );
NAND2_X1 \EXU/_1768_ ( .A1(\EXU/_1131_ ), .A2(\EXU/_0533_ ), .ZN(\EXU/_1140_ ) );
NAND2_X1 \EXU/_1769_ ( .A1(\EXU/_1139_ ), .A2(\EXU/_1140_ ), .ZN(\EXU/_0355_ ) );
NAND2_X1 \EXU/_1770_ ( .A1(\EXU/_1127_ ), .A2(\EXU/_0402_ ), .ZN(\EXU/_1141_ ) );
NAND2_X1 \EXU/_1771_ ( .A1(\EXU/_1131_ ), .A2(\EXU/_0534_ ), .ZN(\EXU/_1142_ ) );
NAND2_X1 \EXU/_1772_ ( .A1(\EXU/_1141_ ), .A2(\EXU/_1142_ ), .ZN(\EXU/_0356_ ) );
NAND2_X1 \EXU/_1773_ ( .A1(\EXU/_1127_ ), .A2(\EXU/_0403_ ), .ZN(\EXU/_1143_ ) );
NAND2_X1 \EXU/_1774_ ( .A1(\EXU/_1131_ ), .A2(\EXU/_0535_ ), .ZN(\EXU/_1144_ ) );
NAND2_X1 \EXU/_1775_ ( .A1(\EXU/_1143_ ), .A2(\EXU/_1144_ ), .ZN(\EXU/_0357_ ) );
NAND2_X1 \EXU/_1776_ ( .A1(\EXU/_1127_ ), .A2(\EXU/_0404_ ), .ZN(\EXU/_1145_ ) );
NAND2_X1 \EXU/_1777_ ( .A1(\EXU/_1131_ ), .A2(\EXU/_0536_ ), .ZN(\EXU/_1146_ ) );
NAND2_X1 \EXU/_1778_ ( .A1(\EXU/_1145_ ), .A2(\EXU/_1146_ ), .ZN(\EXU/_0358_ ) );
NAND2_X1 \EXU/_1779_ ( .A1(\EXU/_1127_ ), .A2(\EXU/_0405_ ), .ZN(\EXU/_1147_ ) );
NAND2_X1 \EXU/_1780_ ( .A1(\EXU/_1131_ ), .A2(\EXU/_0537_ ), .ZN(\EXU/_1148_ ) );
NAND2_X1 \EXU/_1781_ ( .A1(\EXU/_1147_ ), .A2(\EXU/_1148_ ), .ZN(\EXU/_0359_ ) );
BUF_X4 \EXU/_1782_ ( .A(\EXU/_1103_ ), .Z(\EXU/_1149_ ) );
NAND2_X1 \EXU/_1783_ ( .A1(\EXU/_1149_ ), .A2(\EXU/_0407_ ), .ZN(\EXU/_1150_ ) );
NAND2_X1 \EXU/_1784_ ( .A1(\EXU/_1131_ ), .A2(\EXU/_0539_ ), .ZN(\EXU/_1151_ ) );
NAND2_X1 \EXU/_1785_ ( .A1(\EXU/_1150_ ), .A2(\EXU/_1151_ ), .ZN(\EXU/_0361_ ) );
NAND2_X1 \EXU/_1786_ ( .A1(\EXU/_1149_ ), .A2(\EXU/_0408_ ), .ZN(\EXU/_1152_ ) );
BUF_X4 \EXU/_1787_ ( .A(\EXU/_1106_ ), .Z(\EXU/_1153_ ) );
NAND2_X1 \EXU/_1788_ ( .A1(\EXU/_1153_ ), .A2(\EXU/_0540_ ), .ZN(\EXU/_1154_ ) );
NAND2_X1 \EXU/_1789_ ( .A1(\EXU/_1152_ ), .A2(\EXU/_1154_ ), .ZN(\EXU/_0362_ ) );
NAND2_X1 \EXU/_1790_ ( .A1(\EXU/_1149_ ), .A2(\EXU/_0409_ ), .ZN(\EXU/_1155_ ) );
NAND2_X1 \EXU/_1791_ ( .A1(\EXU/_1153_ ), .A2(\EXU/_0541_ ), .ZN(\EXU/_1156_ ) );
NAND2_X1 \EXU/_1792_ ( .A1(\EXU/_1155_ ), .A2(\EXU/_1156_ ), .ZN(\EXU/_0363_ ) );
NAND2_X1 \EXU/_1793_ ( .A1(\EXU/_1149_ ), .A2(\EXU/_0410_ ), .ZN(\EXU/_1157_ ) );
NAND2_X1 \EXU/_1794_ ( .A1(\EXU/_1153_ ), .A2(\EXU/_0542_ ), .ZN(\EXU/_1158_ ) );
NAND2_X1 \EXU/_1795_ ( .A1(\EXU/_1157_ ), .A2(\EXU/_1158_ ), .ZN(\EXU/_0364_ ) );
NAND2_X1 \EXU/_1796_ ( .A1(\EXU/_1149_ ), .A2(\EXU/_0411_ ), .ZN(\EXU/_1159_ ) );
NAND2_X1 \EXU/_1797_ ( .A1(\EXU/_1153_ ), .A2(\EXU/_0543_ ), .ZN(\EXU/_1160_ ) );
NAND2_X1 \EXU/_1798_ ( .A1(\EXU/_1159_ ), .A2(\EXU/_1160_ ), .ZN(\EXU/_0365_ ) );
NAND2_X1 \EXU/_1799_ ( .A1(\EXU/_1149_ ), .A2(\EXU/_0412_ ), .ZN(\EXU/_1161_ ) );
NAND2_X1 \EXU/_1800_ ( .A1(\EXU/_1153_ ), .A2(\EXU/_0544_ ), .ZN(\EXU/_1162_ ) );
NAND2_X1 \EXU/_1801_ ( .A1(\EXU/_1161_ ), .A2(\EXU/_1162_ ), .ZN(\EXU/_0366_ ) );
NAND2_X1 \EXU/_1802_ ( .A1(\EXU/_1149_ ), .A2(\EXU/_0413_ ), .ZN(\EXU/_1163_ ) );
NAND2_X1 \EXU/_1803_ ( .A1(\EXU/_1153_ ), .A2(\EXU/_0545_ ), .ZN(\EXU/_1164_ ) );
NAND2_X1 \EXU/_1804_ ( .A1(\EXU/_1163_ ), .A2(\EXU/_1164_ ), .ZN(\EXU/_0367_ ) );
NAND2_X1 \EXU/_1805_ ( .A1(\EXU/_1149_ ), .A2(\EXU/_0414_ ), .ZN(\EXU/_1165_ ) );
NAND2_X1 \EXU/_1806_ ( .A1(\EXU/_1153_ ), .A2(\EXU/_0546_ ), .ZN(\EXU/_1166_ ) );
NAND2_X1 \EXU/_1807_ ( .A1(\EXU/_1165_ ), .A2(\EXU/_1166_ ), .ZN(\EXU/_0368_ ) );
NAND2_X1 \EXU/_1808_ ( .A1(\EXU/_1106_ ), .A2(\EXU/_0547_ ), .ZN(\EXU/_1167_ ) );
INV_X1 \EXU/_1809_ ( .A(\EXU/_1103_ ), .ZN(\EXU/_1168_ ) );
INV_X1 \EXU/_1810_ ( .A(\EXU/_0415_ ), .ZN(\EXU/_1169_ ) );
OAI21_X1 \EXU/_1811_ ( .A(\EXU/_1167_ ), .B1(\EXU/_1168_ ), .B2(\EXU/_1169_ ), .ZN(\EXU/_0369_ ) );
NAND2_X1 \EXU/_1812_ ( .A1(\EXU/_1149_ ), .A2(\EXU/_0416_ ), .ZN(\EXU/_1170_ ) );
NAND2_X1 \EXU/_1813_ ( .A1(\EXU/_1153_ ), .A2(\EXU/_0548_ ), .ZN(\EXU/_1171_ ) );
NAND2_X1 \EXU/_1814_ ( .A1(\EXU/_1170_ ), .A2(\EXU/_1171_ ), .ZN(\EXU/_0370_ ) );
NAND2_X1 \EXU/_1815_ ( .A1(\EXU/_1149_ ), .A2(\EXU/_0418_ ), .ZN(\EXU/_1172_ ) );
NAND2_X1 \EXU/_1816_ ( .A1(\EXU/_1153_ ), .A2(\EXU/_0550_ ), .ZN(\EXU/_1173_ ) );
NAND2_X1 \EXU/_1817_ ( .A1(\EXU/_1172_ ), .A2(\EXU/_1173_ ), .ZN(\EXU/_0372_ ) );
NAND2_X1 \EXU/_1818_ ( .A1(\EXU/_1103_ ), .A2(\EXU/_0419_ ), .ZN(\EXU/_1174_ ) );
NAND2_X1 \EXU/_1819_ ( .A1(\EXU/_1153_ ), .A2(\EXU/_0551_ ), .ZN(\EXU/_1175_ ) );
NAND2_X1 \EXU/_1820_ ( .A1(\EXU/_1174_ ), .A2(\EXU/_1175_ ), .ZN(\EXU/_0373_ ) );
INV_X32 \EXU/_1821_ ( .A(fanout_net_9 ), .ZN(\EXU/_1176_ ) );
NAND2_X1 \EXU/_1822_ ( .A1(\EXU/_1176_ ), .A2(\EXU/_0470_ ), .ZN(\EXU/_1177_ ) );
NAND2_X1 \EXU/_1823_ ( .A1(\EXU/_0438_ ), .A2(fanout_net_9 ), .ZN(\EXU/_1178_ ) );
NAND2_X1 \EXU/_1824_ ( .A1(\EXU/_1177_ ), .A2(\EXU/_1178_ ), .ZN(\EXU/_1179_ ) );
AND2_X1 \EXU/_1825_ ( .A1(\EXU/_0406_ ), .A2(fanout_net_8 ), .ZN(\EXU/_1180_ ) );
INV_X1 \EXU/_1826_ ( .A(\EXU/_1180_ ), .ZN(\EXU/_1181_ ) );
XNOR2_X1 \EXU/_1827_ ( .A(\EXU/_1179_ ), .B(\EXU/_1181_ ), .ZN(\EXU/_1182_ ) );
NAND2_X1 \EXU/_1828_ ( .A1(\EXU/_1176_ ), .A2(\EXU/_0459_ ), .ZN(\EXU/_1183_ ) );
NAND2_X1 \EXU/_1829_ ( .A1(\EXU/_0427_ ), .A2(fanout_net_9 ), .ZN(\EXU/_1184_ ) );
NAND2_X1 \EXU/_1830_ ( .A1(\EXU/_1183_ ), .A2(\EXU/_1184_ ), .ZN(\EXU/_1185_ ) );
AND2_X1 \EXU/_1831_ ( .A1(\EXU/_0395_ ), .A2(fanout_net_8 ), .ZN(\EXU/_1186_ ) );
AND2_X1 \EXU/_1832_ ( .A1(\EXU/_1185_ ), .A2(\EXU/_1186_ ), .ZN(\EXU/_1187_ ) );
XOR2_X1 \EXU/_1833_ ( .A(\EXU/_1182_ ), .B(\EXU/_1187_ ), .Z(\EXU/_0820_ ) );
AND2_X1 \EXU/_1834_ ( .A1(\EXU/_1182_ ), .A2(\EXU/_1187_ ), .ZN(\EXU/_1188_ ) );
AOI21_X1 \EXU/_1835_ ( .A(\EXU/_1181_ ), .B1(\EXU/_1177_ ), .B2(\EXU/_1178_ ), .ZN(\EXU/_1189_ ) );
NOR2_X1 \EXU/_1836_ ( .A1(\EXU/_1188_ ), .A2(\EXU/_1189_ ), .ZN(\EXU/_1190_ ) );
MUX2_X1 \EXU/_1837_ ( .A(\EXU/_0481_ ), .B(\EXU/_0449_ ), .S(fanout_net_9 ), .Z(\EXU/_1191_ ) );
NAND2_X1 \EXU/_1838_ ( .A1(\EXU/_1112_ ), .A2(fanout_net_8 ), .ZN(\EXU/_1192_ ) );
XOR2_X2 \EXU/_1839_ ( .A(\EXU/_1191_ ), .B(\EXU/_1192_ ), .Z(\EXU/_1193_ ) );
XNOR2_X1 \EXU/_1840_ ( .A(\EXU/_1190_ ), .B(\EXU/_1193_ ), .ZN(\EXU/_0831_ ) );
OAI21_X1 \EXU/_1841_ ( .A(\EXU/_1193_ ), .B1(\EXU/_1188_ ), .B2(\EXU/_1189_ ), .ZN(\EXU/_1194_ ) );
NAND2_X1 \EXU/_1842_ ( .A1(\EXU/_1191_ ), .A2(\EXU/_1192_ ), .ZN(\EXU/_1195_ ) );
NAND2_X1 \EXU/_1843_ ( .A1(\EXU/_1194_ ), .A2(\EXU/_1195_ ), .ZN(\EXU/_1196_ ) );
MUX2_X1 \EXU/_1844_ ( .A(\EXU/_0484_ ), .B(\EXU/_0452_ ), .S(fanout_net_9 ), .Z(\EXU/_1197_ ) );
AND2_X1 \EXU/_1845_ ( .A1(\EXU/_0420_ ), .A2(fanout_net_8 ), .ZN(\EXU/_1198_ ) );
XNOR2_X1 \EXU/_1846_ ( .A(\EXU/_1197_ ), .B(\EXU/_1198_ ), .ZN(\EXU/_1199_ ) );
XNOR2_X1 \EXU/_1847_ ( .A(\EXU/_1196_ ), .B(\EXU/_1199_ ), .ZN(\EXU/_0834_ ) );
INV_X1 \EXU/_1848_ ( .A(\EXU/_1193_ ), .ZN(\EXU/_1200_ ) );
NOR3_X1 \EXU/_1849_ ( .A1(\EXU/_1190_ ), .A2(\EXU/_1200_ ), .A3(\EXU/_1199_ ), .ZN(\EXU/_1201_ ) );
NAND2_X1 \EXU/_1850_ ( .A1(\EXU/_1197_ ), .A2(\EXU/_1198_ ), .ZN(\EXU/_1202_ ) );
OAI21_X1 \EXU/_1851_ ( .A(\EXU/_1202_ ), .B1(\EXU/_1199_ ), .B2(\EXU/_1195_ ), .ZN(\EXU/_1203_ ) );
NOR2_X1 \EXU/_1852_ ( .A1(\EXU/_1201_ ), .A2(\EXU/_1203_ ), .ZN(\EXU/_1204_ ) );
MUX2_X1 \EXU/_1853_ ( .A(\EXU/_0485_ ), .B(\EXU/_0453_ ), .S(fanout_net_9 ), .Z(\EXU/_1205_ ) );
AND2_X1 \EXU/_1854_ ( .A1(\EXU/_0421_ ), .A2(fanout_net_8 ), .ZN(\EXU/_1206_ ) );
XOR2_X1 \EXU/_1855_ ( .A(\EXU/_1205_ ), .B(\EXU/_1206_ ), .Z(\EXU/_1207_ ) );
XNOR2_X1 \EXU/_1856_ ( .A(\EXU/_1204_ ), .B(\EXU/_1207_ ), .ZN(\EXU/_0835_ ) );
INV_X1 \EXU/_1857_ ( .A(\EXU/_1204_ ), .ZN(\EXU/_1208_ ) );
AND2_X1 \EXU/_1858_ ( .A1(\EXU/_1208_ ), .A2(\EXU/_1207_ ), .ZN(\EXU/_1209_ ) );
AND2_X1 \EXU/_1859_ ( .A1(\EXU/_1205_ ), .A2(\EXU/_1206_ ), .ZN(\EXU/_1210_ ) );
NOR2_X1 \EXU/_1860_ ( .A1(\EXU/_1209_ ), .A2(\EXU/_1210_ ), .ZN(\EXU/_1211_ ) );
MUX2_X1 \EXU/_1861_ ( .A(\EXU/_0486_ ), .B(\EXU/_0454_ ), .S(fanout_net_9 ), .Z(\EXU/_1212_ ) );
AND2_X1 \EXU/_1862_ ( .A1(\EXU/_0422_ ), .A2(fanout_net_8 ), .ZN(\EXU/_1213_ ) );
XOR2_X2 \EXU/_1863_ ( .A(\EXU/_1212_ ), .B(\EXU/_1213_ ), .Z(\EXU/_0843_ ) );
XNOR2_X1 \EXU/_1864_ ( .A(\EXU/_1211_ ), .B(\EXU/_0843_ ), .ZN(\EXU/_0836_ ) );
AND3_X1 \EXU/_1865_ ( .A1(\EXU/_1208_ ), .A2(\EXU/_1207_ ), .A3(\EXU/_0843_ ), .ZN(\EXU/_0844_ ) );
AND2_X2 \EXU/_1866_ ( .A1(\EXU/_0843_ ), .A2(\EXU/_1210_ ), .ZN(\EXU/_0845_ ) );
AOI21_X1 \EXU/_1867_ ( .A(\EXU/_0845_ ), .B1(\EXU/_1213_ ), .B2(\EXU/_1212_ ), .ZN(\EXU/_0846_ ) );
INV_X1 \EXU/_1868_ ( .A(\EXU/_0846_ ), .ZN(\EXU/_0847_ ) );
NOR2_X1 \EXU/_1869_ ( .A1(\EXU/_0844_ ), .A2(\EXU/_0847_ ), .ZN(\EXU/_0848_ ) );
MUX2_X1 \EXU/_1870_ ( .A(\EXU/_0487_ ), .B(\EXU/_0455_ ), .S(fanout_net_9 ), .Z(\EXU/_0849_ ) );
AND2_X1 \EXU/_1871_ ( .A1(\EXU/_0423_ ), .A2(fanout_net_8 ), .ZN(\EXU/_0850_ ) );
XOR2_X1 \EXU/_1872_ ( .A(\EXU/_0849_ ), .B(\EXU/_0850_ ), .Z(\EXU/_0851_ ) );
XNOR2_X1 \EXU/_1873_ ( .A(\EXU/_0848_ ), .B(\EXU/_0851_ ), .ZN(\EXU/_0837_ ) );
OAI21_X1 \EXU/_1874_ ( .A(\EXU/_0851_ ), .B1(\EXU/_0844_ ), .B2(\EXU/_0847_ ), .ZN(\EXU/_0852_ ) );
NAND2_X1 \EXU/_1875_ ( .A1(\EXU/_0849_ ), .A2(\EXU/_0850_ ), .ZN(\EXU/_0853_ ) );
NAND2_X1 \EXU/_1876_ ( .A1(\EXU/_0852_ ), .A2(\EXU/_0853_ ), .ZN(\EXU/_0854_ ) );
MUX2_X1 \EXU/_1877_ ( .A(\EXU/_0488_ ), .B(\EXU/_0456_ ), .S(fanout_net_9 ), .Z(\EXU/_0855_ ) );
AND2_X1 \EXU/_1878_ ( .A1(\EXU/_0424_ ), .A2(fanout_net_8 ), .ZN(\EXU/_0856_ ) );
XOR2_X1 \EXU/_1879_ ( .A(\EXU/_0855_ ), .B(\EXU/_0856_ ), .Z(\EXU/_0857_ ) );
INV_X1 \EXU/_1880_ ( .A(\EXU/_0857_ ), .ZN(\EXU/_0858_ ) );
XNOR2_X1 \EXU/_1881_ ( .A(\EXU/_0854_ ), .B(\EXU/_0858_ ), .ZN(\EXU/_0838_ ) );
AND2_X1 \EXU/_1882_ ( .A1(\EXU/_0857_ ), .A2(\EXU/_0851_ ), .ZN(\EXU/_0859_ ) );
AND2_X2 \EXU/_1883_ ( .A1(\EXU/_0847_ ), .A2(\EXU/_0859_ ), .ZN(\EXU/_0860_ ) );
AND2_X1 \EXU/_1884_ ( .A1(\EXU/_0855_ ), .A2(\EXU/_0856_ ), .ZN(\EXU/_0861_ ) );
AND3_X1 \EXU/_1885_ ( .A1(\EXU/_0857_ ), .A2(\EXU/_0850_ ), .A3(\EXU/_0849_ ), .ZN(\EXU/_0862_ ) );
OR3_X4 \EXU/_1886_ ( .A1(\EXU/_0860_ ), .A2(\EXU/_0861_ ), .A3(\EXU/_0862_ ), .ZN(\EXU/_0863_ ) );
AND4_X4 \EXU/_1887_ ( .A1(\EXU/_1208_ ), .A2(\EXU/_1207_ ), .A3(\EXU/_0843_ ), .A4(\EXU/_0859_ ), .ZN(\EXU/_0864_ ) );
NOR2_X4 \EXU/_1888_ ( .A1(\EXU/_0863_ ), .A2(\EXU/_0864_ ), .ZN(\EXU/_0865_ ) );
MUX2_X1 \EXU/_1889_ ( .A(\EXU/_0489_ ), .B(\EXU/_0457_ ), .S(fanout_net_9 ), .Z(\EXU/_0866_ ) );
AND2_X1 \EXU/_1890_ ( .A1(\EXU/_0425_ ), .A2(fanout_net_8 ), .ZN(\EXU/_0867_ ) );
XOR2_X1 \EXU/_1891_ ( .A(\EXU/_0866_ ), .B(\EXU/_0867_ ), .Z(\EXU/_0868_ ) );
XNOR2_X1 \EXU/_1892_ ( .A(\EXU/_0865_ ), .B(\EXU/_0868_ ), .ZN(\EXU/_0839_ ) );
INV_X1 \EXU/_1893_ ( .A(\EXU/_0865_ ), .ZN(\EXU/_0869_ ) );
AND2_X1 \EXU/_1894_ ( .A1(\EXU/_0869_ ), .A2(\EXU/_0868_ ), .ZN(\EXU/_0870_ ) );
AND2_X1 \EXU/_1895_ ( .A1(\EXU/_0866_ ), .A2(\EXU/_0867_ ), .ZN(\EXU/_0871_ ) );
NOR2_X1 \EXU/_1896_ ( .A1(\EXU/_0870_ ), .A2(\EXU/_0871_ ), .ZN(\EXU/_0872_ ) );
MUX2_X1 \EXU/_1897_ ( .A(\EXU/_0490_ ), .B(\EXU/_0458_ ), .S(fanout_net_9 ), .Z(\EXU/_0873_ ) );
AND2_X1 \EXU/_1898_ ( .A1(\EXU/_0426_ ), .A2(fanout_net_8 ), .ZN(\EXU/_0874_ ) );
XOR2_X1 \EXU/_1899_ ( .A(\EXU/_0873_ ), .B(\EXU/_0874_ ), .Z(\EXU/_0875_ ) );
XNOR2_X1 \EXU/_1900_ ( .A(\EXU/_0872_ ), .B(\EXU/_0875_ ), .ZN(\EXU/_0840_ ) );
AND2_X1 \EXU/_1901_ ( .A1(\EXU/_0868_ ), .A2(\EXU/_0875_ ), .ZN(\EXU/_0876_ ) );
AND2_X1 \EXU/_1902_ ( .A1(\EXU/_0869_ ), .A2(\EXU/_0876_ ), .ZN(\EXU/_0877_ ) );
AND2_X1 \EXU/_1903_ ( .A1(\EXU/_0875_ ), .A2(\EXU/_0871_ ), .ZN(\EXU/_0878_ ) );
AOI21_X1 \EXU/_1904_ ( .A(\EXU/_0878_ ), .B1(\EXU/_0874_ ), .B2(\EXU/_0873_ ), .ZN(\EXU/_0879_ ) );
INV_X1 \EXU/_1905_ ( .A(\EXU/_0879_ ), .ZN(\EXU/_0880_ ) );
NOR2_X1 \EXU/_1906_ ( .A1(\EXU/_0877_ ), .A2(\EXU/_0880_ ), .ZN(\EXU/_0881_ ) );
MUX2_X1 \EXU/_1907_ ( .A(\EXU/_0460_ ), .B(\EXU/_0428_ ), .S(fanout_net_9 ), .Z(\EXU/_0882_ ) );
AND2_X1 \EXU/_1908_ ( .A1(\EXU/_0396_ ), .A2(fanout_net_8 ), .ZN(\EXU/_0883_ ) );
XOR2_X1 \EXU/_1909_ ( .A(\EXU/_0882_ ), .B(\EXU/_0883_ ), .Z(\EXU/_0884_ ) );
XNOR2_X1 \EXU/_1910_ ( .A(\EXU/_0881_ ), .B(\EXU/_0884_ ), .ZN(\EXU/_0810_ ) );
OAI21_X1 \EXU/_1911_ ( .A(\EXU/_0884_ ), .B1(\EXU/_0877_ ), .B2(\EXU/_0880_ ), .ZN(\EXU/_0885_ ) );
AND2_X1 \EXU/_1912_ ( .A1(\EXU/_0882_ ), .A2(\EXU/_0883_ ), .ZN(\EXU/_0886_ ) );
INV_X1 \EXU/_1913_ ( .A(\EXU/_0886_ ), .ZN(\EXU/_0887_ ) );
AND2_X1 \EXU/_1914_ ( .A1(\EXU/_0885_ ), .A2(\EXU/_0887_ ), .ZN(\EXU/_0888_ ) );
MUX2_X1 \EXU/_1915_ ( .A(\EXU/_0461_ ), .B(\EXU/_0429_ ), .S(fanout_net_9 ), .Z(\EXU/_0889_ ) );
AND2_X1 \EXU/_1916_ ( .A1(\EXU/_0397_ ), .A2(fanout_net_8 ), .ZN(\EXU/_0890_ ) );
XOR2_X1 \EXU/_1917_ ( .A(\EXU/_0889_ ), .B(\EXU/_0890_ ), .Z(\EXU/_0891_ ) );
XNOR2_X1 \EXU/_1918_ ( .A(\EXU/_0888_ ), .B(\EXU/_0891_ ), .ZN(\EXU/_0811_ ) );
AND2_X1 \EXU/_1919_ ( .A1(\EXU/_0891_ ), .A2(\EXU/_0884_ ), .ZN(\EXU/_0892_ ) );
AND2_X1 \EXU/_1920_ ( .A1(\EXU/_0876_ ), .A2(\EXU/_0892_ ), .ZN(\EXU/_0893_ ) );
INV_X1 \EXU/_1921_ ( .A(\EXU/_0893_ ), .ZN(\EXU/_0894_ ) );
NOR2_X1 \EXU/_1922_ ( .A1(\EXU/_0865_ ), .A2(\EXU/_0894_ ), .ZN(\EXU/_0895_ ) );
NAND2_X1 \EXU/_1923_ ( .A1(\EXU/_0880_ ), .A2(\EXU/_0892_ ), .ZN(\EXU/_0896_ ) );
AND2_X1 \EXU/_1924_ ( .A1(\EXU/_0891_ ), .A2(\EXU/_0886_ ), .ZN(\EXU/_0897_ ) );
AOI21_X1 \EXU/_1925_ ( .A(\EXU/_0897_ ), .B1(\EXU/_0890_ ), .B2(\EXU/_0889_ ), .ZN(\EXU/_0898_ ) );
AND2_X1 \EXU/_1926_ ( .A1(\EXU/_0896_ ), .A2(\EXU/_0898_ ), .ZN(\EXU/_0899_ ) );
INV_X1 \EXU/_1927_ ( .A(\EXU/_0899_ ), .ZN(\EXU/_0900_ ) );
NOR2_X1 \EXU/_1928_ ( .A1(\EXU/_0895_ ), .A2(\EXU/_0900_ ), .ZN(\EXU/_0901_ ) );
MUX2_X1 \EXU/_1929_ ( .A(\EXU/_0462_ ), .B(\EXU/_0430_ ), .S(fanout_net_9 ), .Z(\EXU/_0902_ ) );
AND2_X1 \EXU/_1930_ ( .A1(\EXU/_0398_ ), .A2(fanout_net_8 ), .ZN(\EXU/_0903_ ) );
XOR2_X1 \EXU/_1931_ ( .A(\EXU/_0902_ ), .B(\EXU/_0903_ ), .Z(\EXU/_0904_ ) );
XNOR2_X1 \EXU/_1932_ ( .A(\EXU/_0901_ ), .B(\EXU/_0904_ ), .ZN(\EXU/_0812_ ) );
OAI21_X1 \EXU/_1933_ ( .A(\EXU/_0904_ ), .B1(\EXU/_0895_ ), .B2(\EXU/_0900_ ), .ZN(\EXU/_0905_ ) );
AND2_X1 \EXU/_1934_ ( .A1(\EXU/_0902_ ), .A2(\EXU/_0903_ ), .ZN(\EXU/_0906_ ) );
INV_X1 \EXU/_1935_ ( .A(\EXU/_0906_ ), .ZN(\EXU/_0907_ ) );
AND2_X1 \EXU/_1936_ ( .A1(\EXU/_0905_ ), .A2(\EXU/_0907_ ), .ZN(\EXU/_0908_ ) );
MUX2_X1 \EXU/_1937_ ( .A(\EXU/_0463_ ), .B(\EXU/_0431_ ), .S(fanout_net_9 ), .Z(\EXU/_0909_ ) );
AND2_X1 \EXU/_1938_ ( .A1(\EXU/_0399_ ), .A2(fanout_net_8 ), .ZN(\EXU/_0910_ ) );
XOR2_X2 \EXU/_1939_ ( .A(\EXU/_0909_ ), .B(\EXU/_0910_ ), .Z(\EXU/_0911_ ) );
XNOR2_X1 \EXU/_1940_ ( .A(\EXU/_0908_ ), .B(\EXU/_0911_ ), .ZN(\EXU/_0813_ ) );
AND2_X1 \EXU/_1941_ ( .A1(\EXU/_0904_ ), .A2(\EXU/_0911_ ), .ZN(\EXU/_0912_ ) );
OAI21_X1 \EXU/_1942_ ( .A(\EXU/_0912_ ), .B1(\EXU/_0895_ ), .B2(\EXU/_0900_ ), .ZN(\EXU/_0913_ ) );
AND2_X2 \EXU/_1943_ ( .A1(\EXU/_0911_ ), .A2(\EXU/_0906_ ), .ZN(\EXU/_0914_ ) );
AOI21_X1 \EXU/_1944_ ( .A(\EXU/_0914_ ), .B1(\EXU/_0910_ ), .B2(\EXU/_0909_ ), .ZN(\EXU/_0915_ ) );
AND2_X1 \EXU/_1945_ ( .A1(\EXU/_0913_ ), .A2(\EXU/_0915_ ), .ZN(\EXU/_0916_ ) );
MUX2_X1 \EXU/_1946_ ( .A(\EXU/_0464_ ), .B(\EXU/_0432_ ), .S(fanout_net_9 ), .Z(\EXU/_0917_ ) );
AND2_X1 \EXU/_1947_ ( .A1(\EXU/_0400_ ), .A2(fanout_net_8 ), .ZN(\EXU/_0918_ ) );
XOR2_X1 \EXU/_1948_ ( .A(\EXU/_0917_ ), .B(\EXU/_0918_ ), .Z(\EXU/_0919_ ) );
XNOR2_X1 \EXU/_1949_ ( .A(\EXU/_0916_ ), .B(\EXU/_0919_ ), .ZN(\EXU/_0814_ ) );
INV_X1 \EXU/_1950_ ( .A(\EXU/_0919_ ), .ZN(\EXU/_0920_ ) );
AOI21_X1 \EXU/_1951_ ( .A(\EXU/_0920_ ), .B1(\EXU/_0913_ ), .B2(\EXU/_0915_ ), .ZN(\EXU/_0921_ ) );
AND2_X1 \EXU/_1952_ ( .A1(\EXU/_0917_ ), .A2(\EXU/_0918_ ), .ZN(\EXU/_0922_ ) );
NOR2_X1 \EXU/_1953_ ( .A1(\EXU/_0921_ ), .A2(\EXU/_0922_ ), .ZN(\EXU/_0923_ ) );
MUX2_X1 \EXU/_1954_ ( .A(\EXU/_0465_ ), .B(\EXU/_0433_ ), .S(fanout_net_9 ), .Z(\EXU/_0924_ ) );
AND2_X1 \EXU/_1955_ ( .A1(\EXU/_0401_ ), .A2(fanout_net_8 ), .ZN(\EXU/_0925_ ) );
XOR2_X1 \EXU/_1956_ ( .A(\EXU/_0924_ ), .B(\EXU/_0925_ ), .Z(\EXU/_0926_ ) );
XNOR2_X1 \EXU/_1957_ ( .A(\EXU/_0923_ ), .B(\EXU/_0926_ ), .ZN(\EXU/_0815_ ) );
NAND3_X1 \EXU/_1958_ ( .A1(\EXU/_0912_ ), .A2(\EXU/_0919_ ), .A3(\EXU/_0926_ ), .ZN(\EXU/_0927_ ) );
NOR3_X4 \EXU/_1959_ ( .A1(\EXU/_0865_ ), .A2(\EXU/_0894_ ), .A3(\EXU/_0927_ ), .ZN(\EXU/_0928_ ) );
AOI21_X1 \EXU/_1960_ ( .A(\EXU/_0927_ ), .B1(\EXU/_0896_ ), .B2(\EXU/_0898_ ), .ZN(\EXU/_0929_ ) );
AND2_X1 \EXU/_1961_ ( .A1(\EXU/_0924_ ), .A2(\EXU/_0925_ ), .ZN(\EXU/_0930_ ) );
INV_X1 \EXU/_1962_ ( .A(\EXU/_0915_ ), .ZN(\EXU/_0931_ ) );
AND3_X2 \EXU/_1963_ ( .A1(\EXU/_0931_ ), .A2(\EXU/_0919_ ), .A3(\EXU/_0926_ ), .ZN(\EXU/_0932_ ) );
AND2_X1 \EXU/_1964_ ( .A1(\EXU/_0926_ ), .A2(\EXU/_0922_ ), .ZN(\EXU/_0933_ ) );
NOR4_X2 \EXU/_1965_ ( .A1(\EXU/_0929_ ), .A2(\EXU/_0930_ ), .A3(\EXU/_0932_ ), .A4(\EXU/_0933_ ), .ZN(\EXU/_0934_ ) );
INV_X1 \EXU/_1966_ ( .A(\EXU/_0934_ ), .ZN(\EXU/_0935_ ) );
NOR2_X4 \EXU/_1967_ ( .A1(\EXU/_0928_ ), .A2(\EXU/_0935_ ), .ZN(\EXU/_0936_ ) );
MUX2_X1 \EXU/_1968_ ( .A(\EXU/_0466_ ), .B(\EXU/_0434_ ), .S(fanout_net_9 ), .Z(\EXU/_0937_ ) );
AND2_X1 \EXU/_1969_ ( .A1(\EXU/_0402_ ), .A2(fanout_net_8 ), .ZN(\EXU/_0938_ ) );
XOR2_X1 \EXU/_1970_ ( .A(\EXU/_0937_ ), .B(\EXU/_0938_ ), .Z(\EXU/_0939_ ) );
XNOR2_X1 \EXU/_1971_ ( .A(\EXU/_0936_ ), .B(\EXU/_0939_ ), .ZN(\EXU/_0816_ ) );
OAI21_X1 \EXU/_1972_ ( .A(\EXU/_0939_ ), .B1(\EXU/_0928_ ), .B2(\EXU/_0935_ ), .ZN(\EXU/_0940_ ) );
NAND2_X1 \EXU/_1973_ ( .A1(\EXU/_0937_ ), .A2(\EXU/_0938_ ), .ZN(\EXU/_0941_ ) );
NAND2_X1 \EXU/_1974_ ( .A1(\EXU/_0940_ ), .A2(\EXU/_0941_ ), .ZN(\EXU/_0942_ ) );
NAND2_X1 \EXU/_1975_ ( .A1(\EXU/_1176_ ), .A2(\EXU/_0467_ ), .ZN(\EXU/_0943_ ) );
NAND2_X1 \EXU/_1976_ ( .A1(\EXU/_0435_ ), .A2(fanout_net_9 ), .ZN(\EXU/_0944_ ) );
NAND2_X1 \EXU/_1977_ ( .A1(\EXU/_0943_ ), .A2(\EXU/_0944_ ), .ZN(\EXU/_0945_ ) );
AND2_X1 \EXU/_1978_ ( .A1(\EXU/_0403_ ), .A2(fanout_net_8 ), .ZN(\EXU/_0946_ ) );
XOR2_X1 \EXU/_1979_ ( .A(\EXU/_0945_ ), .B(\EXU/_0946_ ), .Z(\EXU/_0947_ ) );
INV_X1 \EXU/_1980_ ( .A(\EXU/_0947_ ), .ZN(\EXU/_0948_ ) );
XNOR2_X1 \EXU/_1981_ ( .A(\EXU/_0942_ ), .B(\EXU/_0948_ ), .ZN(\EXU/_0817_ ) );
NOR2_X1 \EXU/_1982_ ( .A1(\EXU/_0940_ ), .A2(\EXU/_0948_ ), .ZN(\EXU/_0949_ ) );
AND3_X1 \EXU/_1983_ ( .A1(\EXU/_0947_ ), .A2(\EXU/_0938_ ), .A3(\EXU/_0937_ ), .ZN(\EXU/_0950_ ) );
AND2_X1 \EXU/_1984_ ( .A1(\EXU/_0945_ ), .A2(\EXU/_0946_ ), .ZN(\EXU/_0951_ ) );
OR2_X1 \EXU/_1985_ ( .A1(\EXU/_0950_ ), .A2(\EXU/_0951_ ), .ZN(\EXU/_0952_ ) );
NOR2_X1 \EXU/_1986_ ( .A1(\EXU/_0949_ ), .A2(\EXU/_0952_ ), .ZN(\EXU/_0953_ ) );
MUX2_X1 \EXU/_1987_ ( .A(\EXU/_0468_ ), .B(\EXU/_0436_ ), .S(fanout_net_9 ), .Z(\EXU/_0954_ ) );
AND2_X1 \EXU/_1988_ ( .A1(\EXU/_0404_ ), .A2(fanout_net_8 ), .ZN(\EXU/_0955_ ) );
XOR2_X1 \EXU/_1989_ ( .A(\EXU/_0954_ ), .B(\EXU/_0955_ ), .Z(\EXU/_0956_ ) );
XNOR2_X1 \EXU/_1990_ ( .A(\EXU/_0953_ ), .B(\EXU/_0956_ ), .ZN(\EXU/_0818_ ) );
OAI21_X1 \EXU/_1991_ ( .A(\EXU/_0956_ ), .B1(\EXU/_0949_ ), .B2(\EXU/_0952_ ), .ZN(\EXU/_0957_ ) );
NAND2_X1 \EXU/_1992_ ( .A1(\EXU/_0954_ ), .A2(\EXU/_0955_ ), .ZN(\EXU/_0958_ ) );
NAND2_X1 \EXU/_1993_ ( .A1(\EXU/_0957_ ), .A2(\EXU/_0958_ ), .ZN(\EXU/_0959_ ) );
MUX2_X1 \EXU/_1994_ ( .A(\EXU/_0469_ ), .B(\EXU/_0437_ ), .S(fanout_net_9 ), .Z(\EXU/_0960_ ) );
AND2_X1 \EXU/_1995_ ( .A1(\EXU/_0405_ ), .A2(fanout_net_8 ), .ZN(\EXU/_0961_ ) );
XOR2_X1 \EXU/_1996_ ( .A(\EXU/_0960_ ), .B(\EXU/_0961_ ), .Z(\EXU/_0962_ ) );
INV_X1 \EXU/_1997_ ( .A(\EXU/_0962_ ), .ZN(\EXU/_0963_ ) );
XNOR2_X1 \EXU/_1998_ ( .A(\EXU/_0959_ ), .B(\EXU/_0963_ ), .ZN(\EXU/_0819_ ) );
AND2_X1 \EXU/_1999_ ( .A1(\EXU/_0956_ ), .A2(\EXU/_0962_ ), .ZN(\EXU/_0964_ ) );
NAND3_X1 \EXU/_2000_ ( .A1(\EXU/_0964_ ), .A2(\EXU/_0939_ ), .A3(\EXU/_0947_ ), .ZN(\EXU/_0965_ ) );
OR2_X1 \EXU/_2001_ ( .A1(\EXU/_0936_ ), .A2(\EXU/_0965_ ), .ZN(\EXU/_0966_ ) );
OAI21_X1 \EXU/_2002_ ( .A(\EXU/_0964_ ), .B1(\EXU/_0950_ ), .B2(\EXU/_0951_ ), .ZN(\EXU/_0967_ ) );
NAND2_X1 \EXU/_2003_ ( .A1(\EXU/_0960_ ), .A2(\EXU/_0961_ ), .ZN(\EXU/_0968_ ) );
NAND3_X1 \EXU/_2004_ ( .A1(\EXU/_0962_ ), .A2(\EXU/_0955_ ), .A3(\EXU/_0954_ ), .ZN(\EXU/_0969_ ) );
AND3_X1 \EXU/_2005_ ( .A1(\EXU/_0967_ ), .A2(\EXU/_0968_ ), .A3(\EXU/_0969_ ), .ZN(\EXU/_0970_ ) );
NAND2_X1 \EXU/_2006_ ( .A1(\EXU/_0966_ ), .A2(\EXU/_0970_ ), .ZN(\EXU/_0971_ ) );
MUX2_X1 \EXU/_2007_ ( .A(\EXU/_0471_ ), .B(\EXU/_0439_ ), .S(fanout_net_9 ), .Z(\EXU/_0972_ ) );
AND2_X1 \EXU/_2008_ ( .A1(\EXU/_0407_ ), .A2(fanout_net_8 ), .ZN(\EXU/_0973_ ) );
XOR2_X1 \EXU/_2009_ ( .A(\EXU/_0972_ ), .B(\EXU/_0973_ ), .Z(\EXU/_0974_ ) );
INV_X1 \EXU/_2010_ ( .A(\EXU/_0974_ ), .ZN(\EXU/_0975_ ) );
XNOR2_X1 \EXU/_2011_ ( .A(\EXU/_0971_ ), .B(\EXU/_0975_ ), .ZN(\EXU/_0821_ ) );
AOI21_X1 \EXU/_2012_ ( .A(\EXU/_0975_ ), .B1(\EXU/_0966_ ), .B2(\EXU/_0970_ ), .ZN(\EXU/_0976_ ) );
AND2_X1 \EXU/_2013_ ( .A1(\EXU/_0972_ ), .A2(\EXU/_0973_ ), .ZN(\EXU/_0977_ ) );
NOR2_X1 \EXU/_2014_ ( .A1(\EXU/_0976_ ), .A2(\EXU/_0977_ ), .ZN(\EXU/_0978_ ) );
NAND2_X1 \EXU/_2015_ ( .A1(\EXU/_1176_ ), .A2(\EXU/_0472_ ), .ZN(\EXU/_0979_ ) );
NAND2_X1 \EXU/_2016_ ( .A1(\EXU/_0440_ ), .A2(fanout_net_9 ), .ZN(\EXU/_0980_ ) );
NAND2_X1 \EXU/_2017_ ( .A1(\EXU/_0979_ ), .A2(\EXU/_0980_ ), .ZN(\EXU/_0981_ ) );
AND2_X1 \EXU/_2018_ ( .A1(\EXU/_0408_ ), .A2(fanout_net_8 ), .ZN(\EXU/_0982_ ) );
XOR2_X1 \EXU/_2019_ ( .A(\EXU/_0981_ ), .B(\EXU/_0982_ ), .Z(\EXU/_0983_ ) );
XNOR2_X1 \EXU/_2020_ ( .A(\EXU/_0978_ ), .B(\EXU/_0983_ ), .ZN(\EXU/_0822_ ) );
AND3_X1 \EXU/_2021_ ( .A1(\EXU/_0971_ ), .A2(\EXU/_0974_ ), .A3(\EXU/_0983_ ), .ZN(\EXU/_0984_ ) );
AND2_X1 \EXU/_2022_ ( .A1(\EXU/_0983_ ), .A2(\EXU/_0977_ ), .ZN(\EXU/_0985_ ) );
AOI21_X1 \EXU/_2023_ ( .A(\EXU/_0985_ ), .B1(\EXU/_0982_ ), .B2(\EXU/_0981_ ), .ZN(\EXU/_0986_ ) );
INV_X1 \EXU/_2024_ ( .A(\EXU/_0986_ ), .ZN(\EXU/_0987_ ) );
NOR2_X1 \EXU/_2025_ ( .A1(\EXU/_0984_ ), .A2(\EXU/_0987_ ), .ZN(\EXU/_0988_ ) );
MUX2_X1 \EXU/_2026_ ( .A(\EXU/_0473_ ), .B(\EXU/_0441_ ), .S(fanout_net_9 ), .Z(\EXU/_0989_ ) );
AND2_X1 \EXU/_2027_ ( .A1(\EXU/_0409_ ), .A2(fanout_net_8 ), .ZN(\EXU/_0990_ ) );
XOR2_X1 \EXU/_2028_ ( .A(\EXU/_0989_ ), .B(\EXU/_0990_ ), .Z(\EXU/_0991_ ) );
XNOR2_X1 \EXU/_2029_ ( .A(\EXU/_0988_ ), .B(\EXU/_0991_ ), .ZN(\EXU/_0823_ ) );
OAI21_X1 \EXU/_2030_ ( .A(\EXU/_0991_ ), .B1(\EXU/_0984_ ), .B2(\EXU/_0987_ ), .ZN(\EXU/_0992_ ) );
AND2_X1 \EXU/_2031_ ( .A1(\EXU/_0989_ ), .A2(\EXU/_0990_ ), .ZN(\EXU/_0993_ ) );
INV_X1 \EXU/_2032_ ( .A(\EXU/_0993_ ), .ZN(\EXU/_0994_ ) );
NAND2_X1 \EXU/_2033_ ( .A1(\EXU/_0992_ ), .A2(\EXU/_0994_ ), .ZN(\EXU/_0995_ ) );
MUX2_X1 \EXU/_2034_ ( .A(\EXU/_0474_ ), .B(\EXU/_0442_ ), .S(fanout_net_9 ), .Z(\EXU/_0996_ ) );
AND2_X1 \EXU/_2035_ ( .A1(\EXU/_0410_ ), .A2(fanout_net_8 ), .ZN(\EXU/_0997_ ) );
XNOR2_X1 \EXU/_2036_ ( .A(\EXU/_0996_ ), .B(\EXU/_0997_ ), .ZN(\EXU/_0998_ ) );
XNOR2_X1 \EXU/_2037_ ( .A(\EXU/_0995_ ), .B(\EXU/_0998_ ), .ZN(\EXU/_0824_ ) );
NAND2_X1 \EXU/_2038_ ( .A1(\EXU/_0996_ ), .A2(\EXU/_0997_ ), .ZN(\EXU/_0999_ ) );
OR2_X1 \EXU/_2039_ ( .A1(\EXU/_0996_ ), .A2(\EXU/_0997_ ), .ZN(\EXU/_1000_ ) );
AND3_X1 \EXU/_2040_ ( .A1(\EXU/_0991_ ), .A2(\EXU/_0999_ ), .A3(\EXU/_1000_ ), .ZN(\EXU/_1001_ ) );
NAND3_X1 \EXU/_2041_ ( .A1(\EXU/_1001_ ), .A2(\EXU/_0974_ ), .A3(\EXU/_0983_ ), .ZN(\EXU/_1002_ ) );
NOR3_X4 \EXU/_2042_ ( .A1(\EXU/_0936_ ), .A2(\EXU/_0965_ ), .A3(\EXU/_1002_ ), .ZN(\EXU/_1003_ ) );
AOI22_X1 \EXU/_2043_ ( .A1(\EXU/_0987_ ), .A2(\EXU/_1001_ ), .B1(\EXU/_0993_ ), .B2(\EXU/_1000_ ), .ZN(\EXU/_1004_ ) );
OAI211_X2 \EXU/_2044_ ( .A(\EXU/_1004_ ), .B(\EXU/_0999_ ), .C1(\EXU/_0970_ ), .C2(\EXU/_1002_ ), .ZN(\EXU/_1005_ ) );
NOR2_X4 \EXU/_2045_ ( .A1(\EXU/_1003_ ), .A2(\EXU/_1005_ ), .ZN(\EXU/_1006_ ) );
MUX2_X1 \EXU/_2046_ ( .A(\EXU/_0475_ ), .B(\EXU/_0443_ ), .S(fanout_net_9 ), .Z(\EXU/_1007_ ) );
AND2_X1 \EXU/_2047_ ( .A1(\EXU/_0411_ ), .A2(fanout_net_8 ), .ZN(\EXU/_1008_ ) );
XOR2_X1 \EXU/_2048_ ( .A(\EXU/_1007_ ), .B(\EXU/_1008_ ), .Z(\EXU/_1009_ ) );
XNOR2_X1 \EXU/_2049_ ( .A(\EXU/_1006_ ), .B(\EXU/_1009_ ), .ZN(\EXU/_0825_ ) );
OAI21_X1 \EXU/_2050_ ( .A(\EXU/_1009_ ), .B1(\EXU/_1003_ ), .B2(\EXU/_1005_ ), .ZN(\EXU/_1010_ ) );
INV_X1 \EXU/_2051_ ( .A(\EXU/_1010_ ), .ZN(\EXU/_1011_ ) );
AND2_X1 \EXU/_2052_ ( .A1(\EXU/_1007_ ), .A2(\EXU/_1008_ ), .ZN(\EXU/_1012_ ) );
NOR2_X1 \EXU/_2053_ ( .A1(\EXU/_1011_ ), .A2(\EXU/_1012_ ), .ZN(\EXU/_1013_ ) );
MUX2_X1 \EXU/_2054_ ( .A(\EXU/_0476_ ), .B(\EXU/_0444_ ), .S(fanout_net_9 ), .Z(\EXU/_1014_ ) );
AND2_X1 \EXU/_2055_ ( .A1(\EXU/_0412_ ), .A2(fanout_net_8 ), .ZN(\EXU/_1015_ ) );
XOR2_X1 \EXU/_2056_ ( .A(\EXU/_1014_ ), .B(\EXU/_1015_ ), .Z(\EXU/_1016_ ) );
XNOR2_X1 \EXU/_2057_ ( .A(\EXU/_1013_ ), .B(\EXU/_1016_ ), .ZN(\EXU/_0826_ ) );
NAND2_X1 \EXU/_2058_ ( .A1(\EXU/_1016_ ), .A2(\EXU/_1009_ ), .ZN(\EXU/_1017_ ) );
NOR2_X1 \EXU/_2059_ ( .A1(\EXU/_1006_ ), .A2(\EXU/_1017_ ), .ZN(\EXU/_1018_ ) );
AND2_X1 \EXU/_2060_ ( .A1(\EXU/_1014_ ), .A2(\EXU/_1015_ ), .ZN(\EXU/_1019_ ) );
AOI21_X1 \EXU/_2061_ ( .A(\EXU/_1019_ ), .B1(\EXU/_1016_ ), .B2(\EXU/_1012_ ), .ZN(\EXU/_1020_ ) );
INV_X1 \EXU/_2062_ ( .A(\EXU/_1020_ ), .ZN(\EXU/_1021_ ) );
NOR2_X1 \EXU/_2063_ ( .A1(\EXU/_1018_ ), .A2(\EXU/_1021_ ), .ZN(\EXU/_1022_ ) );
MUX2_X1 \EXU/_2064_ ( .A(\EXU/_0477_ ), .B(\EXU/_0445_ ), .S(fanout_net_9 ), .Z(\EXU/_1023_ ) );
AND2_X1 \EXU/_2065_ ( .A1(\EXU/_0413_ ), .A2(fanout_net_8 ), .ZN(\EXU/_1024_ ) );
XOR2_X1 \EXU/_2066_ ( .A(\EXU/_1023_ ), .B(\EXU/_1024_ ), .Z(\EXU/_1025_ ) );
XNOR2_X1 \EXU/_2067_ ( .A(\EXU/_1022_ ), .B(\EXU/_1025_ ), .ZN(\EXU/_0827_ ) );
OAI21_X1 \EXU/_2068_ ( .A(\EXU/_1025_ ), .B1(\EXU/_1018_ ), .B2(\EXU/_1021_ ), .ZN(\EXU/_1026_ ) );
NAND2_X1 \EXU/_2069_ ( .A1(\EXU/_1023_ ), .A2(\EXU/_1024_ ), .ZN(\EXU/_1027_ ) );
NAND2_X1 \EXU/_2070_ ( .A1(\EXU/_1026_ ), .A2(\EXU/_1027_ ), .ZN(\EXU/_1028_ ) );
MUX2_X1 \EXU/_2071_ ( .A(\EXU/_0478_ ), .B(\EXU/_0446_ ), .S(fanout_net_9 ), .Z(\EXU/_1029_ ) );
AND2_X1 \EXU/_2072_ ( .A1(\EXU/_0414_ ), .A2(fanout_net_8 ), .ZN(\EXU/_1030_ ) );
XOR2_X1 \EXU/_2073_ ( .A(\EXU/_1029_ ), .B(\EXU/_1030_ ), .Z(\EXU/_1031_ ) );
INV_X1 \EXU/_2074_ ( .A(\EXU/_1031_ ), .ZN(\EXU/_1032_ ) );
XNOR2_X1 \EXU/_2075_ ( .A(\EXU/_1028_ ), .B(\EXU/_1032_ ), .ZN(\EXU/_0828_ ) );
NAND2_X1 \EXU/_2076_ ( .A1(\EXU/_1031_ ), .A2(\EXU/_1025_ ), .ZN(\EXU/_1033_ ) );
NOR3_X4 \EXU/_2077_ ( .A1(\EXU/_1006_ ), .A2(\EXU/_1017_ ), .A3(\EXU/_1033_ ), .ZN(\EXU/_1034_ ) );
AND2_X1 \EXU/_2078_ ( .A1(\EXU/_1029_ ), .A2(\EXU/_1030_ ), .ZN(\EXU/_1035_ ) );
INV_X1 \EXU/_2079_ ( .A(\EXU/_1035_ ), .ZN(\EXU/_1036_ ) );
OAI221_X1 \EXU/_2080_ ( .A(\EXU/_1036_ ), .B1(\EXU/_1032_ ), .B2(\EXU/_1027_ ), .C1(\EXU/_1020_ ), .C2(\EXU/_1033_ ), .ZN(\EXU/_1037_ ) );
NOR2_X1 \EXU/_2081_ ( .A1(\EXU/_1034_ ), .A2(\EXU/_1037_ ), .ZN(\EXU/_1038_ ) );
NAND2_X1 \EXU/_2082_ ( .A1(\EXU/_0447_ ), .A2(fanout_net_9 ), .ZN(\EXU/_1039_ ) );
INV_X1 \EXU/_2083_ ( .A(\EXU/_0479_ ), .ZN(\EXU/_1040_ ) );
OAI21_X1 \EXU/_2084_ ( .A(\EXU/_1039_ ), .B1(\EXU/_1040_ ), .B2(\EXU/_0068_ ), .ZN(\EXU/_1041_ ) );
AND2_X1 \EXU/_2085_ ( .A1(\EXU/_0415_ ), .A2(fanout_net_8 ), .ZN(\EXU/_1042_ ) );
XOR2_X1 \EXU/_2086_ ( .A(\EXU/_1041_ ), .B(\EXU/_1042_ ), .Z(\EXU/_1043_ ) );
XNOR2_X1 \EXU/_2087_ ( .A(\EXU/_1038_ ), .B(\EXU/_1043_ ), .ZN(\EXU/_0829_ ) );
OAI21_X1 \EXU/_2088_ ( .A(\EXU/_1043_ ), .B1(\EXU/_1034_ ), .B2(\EXU/_1037_ ), .ZN(\EXU/_1044_ ) );
NAND2_X1 \EXU/_2089_ ( .A1(\EXU/_1041_ ), .A2(\EXU/_1042_ ), .ZN(\EXU/_1045_ ) );
NAND2_X1 \EXU/_2090_ ( .A1(\EXU/_1044_ ), .A2(\EXU/_1045_ ), .ZN(\EXU/_1046_ ) );
MUX2_X1 \EXU/_2091_ ( .A(\EXU/_0480_ ), .B(\EXU/_0448_ ), .S(\EXU/_0068_ ), .Z(\EXU/_1047_ ) );
AND2_X1 \EXU/_2092_ ( .A1(\EXU/_0416_ ), .A2(fanout_net_8 ), .ZN(\EXU/_1048_ ) );
XNOR2_X1 \EXU/_2093_ ( .A(\EXU/_1047_ ), .B(\EXU/_1048_ ), .ZN(\EXU/_1049_ ) );
XNOR2_X1 \EXU/_2094_ ( .A(\EXU/_1046_ ), .B(\EXU/_1049_ ), .ZN(\EXU/_0830_ ) );
XOR2_X1 \EXU/_2095_ ( .A(\EXU/_1047_ ), .B(\EXU/_1048_ ), .Z(\EXU/_1050_ ) );
OAI211_X2 \EXU/_2096_ ( .A(\EXU/_1043_ ), .B(\EXU/_1050_ ), .C1(\EXU/_1034_ ), .C2(\EXU/_1037_ ), .ZN(\EXU/_1051_ ) );
NOR2_X1 \EXU/_2097_ ( .A1(\EXU/_1049_ ), .A2(\EXU/_1045_ ), .ZN(\EXU/_1052_ ) );
AOI21_X1 \EXU/_2098_ ( .A(\EXU/_1052_ ), .B1(\EXU/_1048_ ), .B2(\EXU/_1047_ ), .ZN(\EXU/_1053_ ) );
AND2_X2 \EXU/_2099_ ( .A1(\EXU/_1051_ ), .A2(\EXU/_1053_ ), .ZN(\EXU/_1054_ ) );
MUX2_X1 \EXU/_2100_ ( .A(\EXU/_0482_ ), .B(\EXU/_0450_ ), .S(\EXU/_0068_ ), .Z(\EXU/_1055_ ) );
AND2_X1 \EXU/_2101_ ( .A1(\EXU/_0418_ ), .A2(\EXU/_0067_ ), .ZN(\EXU/_1056_ ) );
AND2_X1 \EXU/_2102_ ( .A1(\EXU/_1055_ ), .A2(\EXU/_1056_ ), .ZN(\EXU/_1057_ ) );
NOR2_X1 \EXU/_2103_ ( .A1(\EXU/_1055_ ), .A2(\EXU/_1056_ ), .ZN(\EXU/_1058_ ) );
NOR2_X1 \EXU/_2104_ ( .A1(\EXU/_1057_ ), .A2(\EXU/_1058_ ), .ZN(\EXU/_1059_ ) );
XNOR2_X1 \EXU/_2105_ ( .A(\EXU/_1054_ ), .B(\EXU/_1059_ ), .ZN(\EXU/_0832_ ) );
NOR3_X2 \EXU/_2106_ ( .A1(\EXU/_1054_ ), .A2(\EXU/_1057_ ), .A3(\EXU/_1058_ ), .ZN(\EXU/_1060_ ) );
NOR2_X2 \EXU/_2107_ ( .A1(\EXU/_1060_ ), .A2(\EXU/_1057_ ), .ZN(\EXU/_1061_ ) );
NAND2_X1 \EXU/_2108_ ( .A1(\EXU/_1176_ ), .A2(\EXU/_0483_ ), .ZN(\EXU/_1062_ ) );
NAND2_X1 \EXU/_2109_ ( .A1(\EXU/_0451_ ), .A2(\EXU/_0068_ ), .ZN(\EXU/_1063_ ) );
AND4_X1 \EXU/_2110_ ( .A1(\EXU/_0419_ ), .A2(\EXU/_1062_ ), .A3(\EXU/_0067_ ), .A4(\EXU/_1063_ ), .ZN(\EXU/_1064_ ) );
AOI22_X1 \EXU/_2111_ ( .A1(\EXU/_1062_ ), .A2(\EXU/_1063_ ), .B1(\EXU/_0419_ ), .B2(\EXU/_0067_ ), .ZN(\EXU/_1065_ ) );
OR2_X1 \EXU/_2112_ ( .A1(\EXU/_1064_ ), .A2(\EXU/_1065_ ), .ZN(\EXU/_1066_ ) );
XNOR2_X1 \EXU/_2113_ ( .A(\EXU/_1061_ ), .B(\EXU/_1066_ ), .ZN(\EXU/_0833_ ) );
XOR2_X1 \EXU/_2114_ ( .A(\EXU/_1185_ ), .B(\EXU/_1186_ ), .Z(\EXU/_0809_ ) );
AND2_X1 \EXU/_2115_ ( .A1(\EXU/_0594_ ), .A2(\EXU/_0595_ ), .ZN(\EXU/_1067_ ) );
BUF_X4 \EXU/_2116_ ( .A(\EXU/_1067_ ), .Z(\EXU/_1068_ ) );
BUF_X4 \EXU/_2117_ ( .A(\EXU/_1068_ ), .Z(\EXU/_1069_ ) );
MUX2_X1 \EXU/_2118_ ( .A(\EXU/_0777_ ), .B(\EXU/_0562_ ), .S(\EXU/_1069_ ), .Z(\EXU/_0136_ ) );
MUX2_X1 \EXU/_2119_ ( .A(\EXU/_0788_ ), .B(\EXU/_0573_ ), .S(\EXU/_1069_ ), .Z(\EXU/_0137_ ) );
MUX2_X1 \EXU/_2120_ ( .A(\EXU/_0799_ ), .B(\EXU/_0584_ ), .S(\EXU/_1069_ ), .Z(\EXU/_0138_ ) );
MUX2_X1 \EXU/_2121_ ( .A(\EXU/_0802_ ), .B(\EXU/_0587_ ), .S(\EXU/_1069_ ), .Z(\EXU/_0139_ ) );
MUX2_X1 \EXU/_2122_ ( .A(\EXU/_0803_ ), .B(\EXU/_0588_ ), .S(\EXU/_1069_ ), .Z(\EXU/_0140_ ) );
MUX2_X1 \EXU/_2123_ ( .A(\EXU/_0804_ ), .B(\EXU/_0589_ ), .S(\EXU/_1069_ ), .Z(\EXU/_0141_ ) );
MUX2_X1 \EXU/_2124_ ( .A(\EXU/_0805_ ), .B(\EXU/_0590_ ), .S(\EXU/_1069_ ), .Z(\EXU/_0142_ ) );
MUX2_X1 \EXU/_2125_ ( .A(\EXU/_0806_ ), .B(\EXU/_0591_ ), .S(\EXU/_1069_ ), .Z(\EXU/_0143_ ) );
MUX2_X1 \EXU/_2126_ ( .A(\EXU/_0807_ ), .B(\EXU/_0592_ ), .S(\EXU/_1069_ ), .Z(\EXU/_0144_ ) );
BUF_X4 \EXU/_2127_ ( .A(\EXU/_1068_ ), .Z(\EXU/_1070_ ) );
MUX2_X1 \EXU/_2128_ ( .A(\EXU/_0808_ ), .B(\EXU/_0593_ ), .S(\EXU/_1070_ ), .Z(\EXU/_0145_ ) );
MUX2_X1 \EXU/_2129_ ( .A(\EXU/_0778_ ), .B(\EXU/_0563_ ), .S(\EXU/_1070_ ), .Z(\EXU/_0146_ ) );
MUX2_X1 \EXU/_2130_ ( .A(\EXU/_0779_ ), .B(\EXU/_0564_ ), .S(\EXU/_1070_ ), .Z(\EXU/_0147_ ) );
MUX2_X1 \EXU/_2131_ ( .A(\EXU/_0780_ ), .B(\EXU/_0565_ ), .S(\EXU/_1070_ ), .Z(\EXU/_0148_ ) );
MUX2_X1 \EXU/_2132_ ( .A(\EXU/_0781_ ), .B(\EXU/_0566_ ), .S(\EXU/_1070_ ), .Z(\EXU/_0149_ ) );
MUX2_X1 \EXU/_2133_ ( .A(\EXU/_0782_ ), .B(\EXU/_0567_ ), .S(\EXU/_1070_ ), .Z(\EXU/_0150_ ) );
MUX2_X1 \EXU/_2134_ ( .A(\EXU/_0783_ ), .B(\EXU/_0568_ ), .S(\EXU/_1070_ ), .Z(\EXU/_0151_ ) );
MUX2_X1 \EXU/_2135_ ( .A(\EXU/_0784_ ), .B(\EXU/_0569_ ), .S(\EXU/_1070_ ), .Z(\EXU/_0152_ ) );
MUX2_X1 \EXU/_2136_ ( .A(\EXU/_0785_ ), .B(\EXU/_0570_ ), .S(\EXU/_1070_ ), .Z(\EXU/_0153_ ) );
MUX2_X1 \EXU/_2137_ ( .A(\EXU/_0786_ ), .B(\EXU/_0571_ ), .S(\EXU/_1070_ ), .Z(\EXU/_0154_ ) );
BUF_X4 \EXU/_2138_ ( .A(\EXU/_1068_ ), .Z(\EXU/_1071_ ) );
MUX2_X1 \EXU/_2139_ ( .A(\EXU/_0787_ ), .B(\EXU/_0572_ ), .S(\EXU/_1071_ ), .Z(\EXU/_0155_ ) );
MUX2_X1 \EXU/_2140_ ( .A(\EXU/_0789_ ), .B(\EXU/_0574_ ), .S(\EXU/_1071_ ), .Z(\EXU/_0156_ ) );
MUX2_X1 \EXU/_2141_ ( .A(\EXU/_0790_ ), .B(\EXU/_0575_ ), .S(\EXU/_1071_ ), .Z(\EXU/_0157_ ) );
MUX2_X1 \EXU/_2142_ ( .A(\EXU/_0791_ ), .B(\EXU/_0576_ ), .S(\EXU/_1071_ ), .Z(\EXU/_0158_ ) );
MUX2_X1 \EXU/_2143_ ( .A(\EXU/_0792_ ), .B(\EXU/_0577_ ), .S(\EXU/_1071_ ), .Z(\EXU/_0159_ ) );
MUX2_X1 \EXU/_2144_ ( .A(\EXU/_0793_ ), .B(\EXU/_0578_ ), .S(\EXU/_1071_ ), .Z(\EXU/_0160_ ) );
MUX2_X1 \EXU/_2145_ ( .A(\EXU/_0794_ ), .B(\EXU/_0579_ ), .S(\EXU/_1071_ ), .Z(\EXU/_0161_ ) );
MUX2_X1 \EXU/_2146_ ( .A(\EXU/_0795_ ), .B(\EXU/_0580_ ), .S(\EXU/_1071_ ), .Z(\EXU/_0162_ ) );
MUX2_X1 \EXU/_2147_ ( .A(\EXU/_0796_ ), .B(\EXU/_0581_ ), .S(\EXU/_1071_ ), .Z(\EXU/_0163_ ) );
MUX2_X1 \EXU/_2148_ ( .A(\EXU/_0797_ ), .B(\EXU/_0582_ ), .S(\EXU/_1071_ ), .Z(\EXU/_0164_ ) );
MUX2_X1 \EXU/_2149_ ( .A(\EXU/_0798_ ), .B(\EXU/_0583_ ), .S(\EXU/_1068_ ), .Z(\EXU/_0165_ ) );
MUX2_X1 \EXU/_2150_ ( .A(\EXU/_0800_ ), .B(\EXU/_0585_ ), .S(\EXU/_1068_ ), .Z(\EXU/_0166_ ) );
MUX2_X1 \EXU/_2151_ ( .A(\EXU/_0801_ ), .B(\EXU/_0586_ ), .S(\EXU/_1068_ ), .Z(\EXU/_0167_ ) );
AND2_X1 \EXU/_2152_ ( .A1(\EXU/_0775_ ), .A2(\EXU/_0776_ ), .ZN(\EXU/_1072_ ) );
BUF_X8 \EXU/_2153_ ( .A(\EXU/_1072_ ), .Z(\EXU/_1073_ ) );
BUF_X8 \EXU/_2154_ ( .A(\EXU/_1073_ ), .Z(\EXU/_1074_ ) );
BUF_X4 \EXU/_2155_ ( .A(\EXU/_1074_ ), .Z(\EXU/_1075_ ) );
MUX2_X1 \EXU/_2156_ ( .A(\EXU/_0427_ ), .B(\EXU/_0647_ ), .S(\EXU/_1075_ ), .Z(\EXU/_0170_ ) );
MUX2_X1 \EXU/_2157_ ( .A(\EXU/_0438_ ), .B(\EXU/_0658_ ), .S(\EXU/_1075_ ), .Z(\EXU/_0171_ ) );
MUX2_X1 \EXU/_2158_ ( .A(\EXU/_0449_ ), .B(\EXU/_0669_ ), .S(\EXU/_1075_ ), .Z(\EXU/_0172_ ) );
MUX2_X1 \EXU/_2159_ ( .A(\EXU/_0452_ ), .B(\EXU/_0672_ ), .S(\EXU/_1075_ ), .Z(\EXU/_0173_ ) );
MUX2_X1 \EXU/_2160_ ( .A(\EXU/_0453_ ), .B(\EXU/_0673_ ), .S(\EXU/_1075_ ), .Z(\EXU/_0174_ ) );
MUX2_X1 \EXU/_2161_ ( .A(\EXU/_0454_ ), .B(\EXU/_0674_ ), .S(\EXU/_1075_ ), .Z(\EXU/_0175_ ) );
MUX2_X1 \EXU/_2162_ ( .A(\EXU/_0455_ ), .B(\EXU/_0675_ ), .S(\EXU/_1075_ ), .Z(\EXU/_0176_ ) );
MUX2_X1 \EXU/_2163_ ( .A(\EXU/_0456_ ), .B(\EXU/_0676_ ), .S(\EXU/_1075_ ), .Z(\EXU/_0177_ ) );
MUX2_X1 \EXU/_2164_ ( .A(\EXU/_0457_ ), .B(\EXU/_0677_ ), .S(\EXU/_1075_ ), .Z(\EXU/_0178_ ) );
BUF_X4 \EXU/_2165_ ( .A(\EXU/_1074_ ), .Z(\EXU/_1076_ ) );
MUX2_X1 \EXU/_2166_ ( .A(\EXU/_0458_ ), .B(\EXU/_0678_ ), .S(\EXU/_1076_ ), .Z(\EXU/_0179_ ) );
MUX2_X1 \EXU/_2167_ ( .A(\EXU/_0428_ ), .B(\EXU/_0648_ ), .S(\EXU/_1076_ ), .Z(\EXU/_0180_ ) );
MUX2_X1 \EXU/_2168_ ( .A(\EXU/_0429_ ), .B(\EXU/_0649_ ), .S(\EXU/_1076_ ), .Z(\EXU/_0181_ ) );
MUX2_X1 \EXU/_2169_ ( .A(\EXU/_0430_ ), .B(\EXU/_0650_ ), .S(\EXU/_1076_ ), .Z(\EXU/_0182_ ) );
MUX2_X1 \EXU/_2170_ ( .A(\EXU/_0431_ ), .B(\EXU/_0651_ ), .S(\EXU/_1076_ ), .Z(\EXU/_0183_ ) );
MUX2_X1 \EXU/_2171_ ( .A(\EXU/_0432_ ), .B(\EXU/_0652_ ), .S(\EXU/_1076_ ), .Z(\EXU/_0184_ ) );
MUX2_X1 \EXU/_2172_ ( .A(\EXU/_0433_ ), .B(\EXU/_0653_ ), .S(\EXU/_1076_ ), .Z(\EXU/_0185_ ) );
MUX2_X1 \EXU/_2173_ ( .A(\EXU/_0434_ ), .B(\EXU/_0654_ ), .S(\EXU/_1076_ ), .Z(\EXU/_0186_ ) );
MUX2_X1 \EXU/_2174_ ( .A(\EXU/_0435_ ), .B(\EXU/_0655_ ), .S(\EXU/_1076_ ), .Z(\EXU/_0187_ ) );
MUX2_X1 \EXU/_2175_ ( .A(\EXU/_0436_ ), .B(\EXU/_0656_ ), .S(\EXU/_1076_ ), .Z(\EXU/_0188_ ) );
BUF_X4 \EXU/_2176_ ( .A(\EXU/_1074_ ), .Z(\EXU/_1077_ ) );
MUX2_X1 \EXU/_2177_ ( .A(\EXU/_0437_ ), .B(\EXU/_0657_ ), .S(\EXU/_1077_ ), .Z(\EXU/_0189_ ) );
MUX2_X1 \EXU/_2178_ ( .A(\EXU/_0439_ ), .B(\EXU/_0659_ ), .S(\EXU/_1077_ ), .Z(\EXU/_0190_ ) );
MUX2_X1 \EXU/_2179_ ( .A(\EXU/_0440_ ), .B(\EXU/_0660_ ), .S(\EXU/_1077_ ), .Z(\EXU/_0191_ ) );
MUX2_X1 \EXU/_2180_ ( .A(\EXU/_0441_ ), .B(\EXU/_0661_ ), .S(\EXU/_1077_ ), .Z(\EXU/_0192_ ) );
MUX2_X1 \EXU/_2181_ ( .A(\EXU/_0442_ ), .B(\EXU/_0662_ ), .S(\EXU/_1077_ ), .Z(\EXU/_0193_ ) );
MUX2_X1 \EXU/_2182_ ( .A(\EXU/_0443_ ), .B(\EXU/_0663_ ), .S(\EXU/_1077_ ), .Z(\EXU/_0194_ ) );
MUX2_X1 \EXU/_2183_ ( .A(\EXU/_0444_ ), .B(\EXU/_0664_ ), .S(\EXU/_1077_ ), .Z(\EXU/_0195_ ) );
MUX2_X1 \EXU/_2184_ ( .A(\EXU/_0445_ ), .B(\EXU/_0665_ ), .S(\EXU/_1077_ ), .Z(\EXU/_0196_ ) );
MUX2_X1 \EXU/_2185_ ( .A(\EXU/_0446_ ), .B(\EXU/_0666_ ), .S(\EXU/_1077_ ), .Z(\EXU/_0197_ ) );
MUX2_X1 \EXU/_2186_ ( .A(\EXU/_0447_ ), .B(\EXU/_0667_ ), .S(\EXU/_1077_ ), .Z(\EXU/_0198_ ) );
BUF_X4 \EXU/_2187_ ( .A(\EXU/_1074_ ), .Z(\EXU/_1078_ ) );
MUX2_X1 \EXU/_2188_ ( .A(\EXU/_0448_ ), .B(\EXU/_0668_ ), .S(\EXU/_1078_ ), .Z(\EXU/_0199_ ) );
MUX2_X1 \EXU/_2189_ ( .A(\EXU/_0450_ ), .B(\EXU/_0670_ ), .S(\EXU/_1078_ ), .Z(\EXU/_0200_ ) );
MUX2_X1 \EXU/_2190_ ( .A(\EXU/_0451_ ), .B(\EXU/_0671_ ), .S(\EXU/_1078_ ), .Z(\EXU/_0201_ ) );
MUX2_X1 \EXU/_2191_ ( .A(\EXU/_0459_ ), .B(\EXU/_0679_ ), .S(\EXU/_1078_ ), .Z(\EXU/_0202_ ) );
MUX2_X1 \EXU/_2192_ ( .A(\EXU/_0470_ ), .B(\EXU/_0690_ ), .S(\EXU/_1078_ ), .Z(\EXU/_0203_ ) );
MUX2_X1 \EXU/_2193_ ( .A(\EXU/_0481_ ), .B(\EXU/_0701_ ), .S(\EXU/_1078_ ), .Z(\EXU/_0204_ ) );
MUX2_X1 \EXU/_2194_ ( .A(\EXU/_0484_ ), .B(\EXU/_0704_ ), .S(\EXU/_1078_ ), .Z(\EXU/_0205_ ) );
MUX2_X1 \EXU/_2195_ ( .A(\EXU/_0485_ ), .B(\EXU/_0705_ ), .S(\EXU/_1078_ ), .Z(\EXU/_0206_ ) );
MUX2_X1 \EXU/_2196_ ( .A(\EXU/_0486_ ), .B(\EXU/_0706_ ), .S(\EXU/_1078_ ), .Z(\EXU/_0207_ ) );
MUX2_X1 \EXU/_2197_ ( .A(\EXU/_0487_ ), .B(\EXU/_0707_ ), .S(\EXU/_1078_ ), .Z(\EXU/_0208_ ) );
BUF_X4 \EXU/_2198_ ( .A(\EXU/_1074_ ), .Z(\EXU/_1079_ ) );
MUX2_X1 \EXU/_2199_ ( .A(\EXU/_0488_ ), .B(\EXU/_0708_ ), .S(\EXU/_1079_ ), .Z(\EXU/_0209_ ) );
MUX2_X1 \EXU/_2200_ ( .A(\EXU/_0489_ ), .B(\EXU/_0709_ ), .S(\EXU/_1079_ ), .Z(\EXU/_0210_ ) );
MUX2_X1 \EXU/_2201_ ( .A(\EXU/_0490_ ), .B(\EXU/_0710_ ), .S(\EXU/_1079_ ), .Z(\EXU/_0211_ ) );
MUX2_X1 \EXU/_2202_ ( .A(\EXU/_0460_ ), .B(\EXU/_0680_ ), .S(\EXU/_1079_ ), .Z(\EXU/_0212_ ) );
MUX2_X1 \EXU/_2203_ ( .A(\EXU/_0461_ ), .B(\EXU/_0681_ ), .S(\EXU/_1079_ ), .Z(\EXU/_0213_ ) );
MUX2_X1 \EXU/_2204_ ( .A(\EXU/_0462_ ), .B(\EXU/_0682_ ), .S(\EXU/_1079_ ), .Z(\EXU/_0214_ ) );
MUX2_X1 \EXU/_2205_ ( .A(\EXU/_0463_ ), .B(\EXU/_0683_ ), .S(\EXU/_1079_ ), .Z(\EXU/_0215_ ) );
MUX2_X1 \EXU/_2206_ ( .A(\EXU/_0464_ ), .B(\EXU/_0684_ ), .S(\EXU/_1079_ ), .Z(\EXU/_0216_ ) );
MUX2_X1 \EXU/_2207_ ( .A(\EXU/_0465_ ), .B(\EXU/_0685_ ), .S(\EXU/_1079_ ), .Z(\EXU/_0217_ ) );
MUX2_X1 \EXU/_2208_ ( .A(\EXU/_0466_ ), .B(\EXU/_0686_ ), .S(\EXU/_1079_ ), .Z(\EXU/_0218_ ) );
BUF_X4 \EXU/_2209_ ( .A(\EXU/_1074_ ), .Z(\EXU/_1080_ ) );
MUX2_X1 \EXU/_2210_ ( .A(\EXU/_0467_ ), .B(\EXU/_0687_ ), .S(\EXU/_1080_ ), .Z(\EXU/_0219_ ) );
MUX2_X1 \EXU/_2211_ ( .A(\EXU/_0468_ ), .B(\EXU/_0688_ ), .S(\EXU/_1080_ ), .Z(\EXU/_0220_ ) );
MUX2_X1 \EXU/_2212_ ( .A(\EXU/_0469_ ), .B(\EXU/_0689_ ), .S(\EXU/_1080_ ), .Z(\EXU/_0221_ ) );
MUX2_X1 \EXU/_2213_ ( .A(\EXU/_0471_ ), .B(\EXU/_0691_ ), .S(\EXU/_1080_ ), .Z(\EXU/_0222_ ) );
MUX2_X1 \EXU/_2214_ ( .A(\EXU/_0472_ ), .B(\EXU/_0692_ ), .S(\EXU/_1080_ ), .Z(\EXU/_0223_ ) );
MUX2_X1 \EXU/_2215_ ( .A(\EXU/_0473_ ), .B(\EXU/_0693_ ), .S(\EXU/_1080_ ), .Z(\EXU/_0224_ ) );
MUX2_X1 \EXU/_2216_ ( .A(\EXU/_0474_ ), .B(\EXU/_0694_ ), .S(\EXU/_1080_ ), .Z(\EXU/_0225_ ) );
MUX2_X1 \EXU/_2217_ ( .A(\EXU/_0475_ ), .B(\EXU/_0695_ ), .S(\EXU/_1080_ ), .Z(\EXU/_0226_ ) );
MUX2_X1 \EXU/_2218_ ( .A(\EXU/_0476_ ), .B(\EXU/_0696_ ), .S(\EXU/_1080_ ), .Z(\EXU/_0227_ ) );
MUX2_X1 \EXU/_2219_ ( .A(\EXU/_0477_ ), .B(\EXU/_0697_ ), .S(\EXU/_1080_ ), .Z(\EXU/_0228_ ) );
BUF_X4 \EXU/_2220_ ( .A(\EXU/_1074_ ), .Z(\EXU/_1081_ ) );
MUX2_X1 \EXU/_2221_ ( .A(\EXU/_0478_ ), .B(\EXU/_0698_ ), .S(\EXU/_1081_ ), .Z(\EXU/_0229_ ) );
MUX2_X1 \EXU/_2222_ ( .A(\EXU/_0479_ ), .B(\EXU/_0699_ ), .S(\EXU/_1081_ ), .Z(\EXU/_0230_ ) );
MUX2_X1 \EXU/_2223_ ( .A(\EXU/_0480_ ), .B(\EXU/_0700_ ), .S(\EXU/_1081_ ), .Z(\EXU/_0231_ ) );
MUX2_X1 \EXU/_2224_ ( .A(\EXU/_0482_ ), .B(\EXU/_0702_ ), .S(\EXU/_1081_ ), .Z(\EXU/_0232_ ) );
MUX2_X1 \EXU/_2225_ ( .A(\EXU/_0483_ ), .B(\EXU/_0703_ ), .S(\EXU/_1081_ ), .Z(\EXU/_0233_ ) );
MUX2_X1 \EXU/_2226_ ( .A(\EXU/_0527_ ), .B(\EXU/_0711_ ), .S(\EXU/_1081_ ), .Z(\EXU/_0234_ ) );
MUX2_X1 \EXU/_2227_ ( .A(\EXU/_0538_ ), .B(\EXU/_0722_ ), .S(\EXU/_1081_ ), .Z(\EXU/_0235_ ) );
MUX2_X1 \EXU/_2228_ ( .A(\EXU/_0549_ ), .B(\EXU/_0733_ ), .S(\EXU/_1081_ ), .Z(\EXU/_0236_ ) );
MUX2_X1 \EXU/_2229_ ( .A(\EXU/_0552_ ), .B(\EXU/_0736_ ), .S(\EXU/_1081_ ), .Z(\EXU/_0237_ ) );
MUX2_X1 \EXU/_2230_ ( .A(\EXU/_0553_ ), .B(\EXU/_0737_ ), .S(\EXU/_1081_ ), .Z(\EXU/_0238_ ) );
BUF_X4 \EXU/_2231_ ( .A(\EXU/_1074_ ), .Z(\EXU/_1082_ ) );
MUX2_X1 \EXU/_2232_ ( .A(\EXU/_0554_ ), .B(\EXU/_0738_ ), .S(\EXU/_1082_ ), .Z(\EXU/_0239_ ) );
MUX2_X1 \EXU/_2233_ ( .A(\EXU/_0555_ ), .B(\EXU/_0739_ ), .S(\EXU/_1082_ ), .Z(\EXU/_0240_ ) );
MUX2_X1 \EXU/_2234_ ( .A(\EXU/_0556_ ), .B(\EXU/_0740_ ), .S(\EXU/_1082_ ), .Z(\EXU/_0241_ ) );
MUX2_X1 \EXU/_2235_ ( .A(\EXU/_0557_ ), .B(\EXU/_0741_ ), .S(\EXU/_1082_ ), .Z(\EXU/_0242_ ) );
MUX2_X1 \EXU/_2236_ ( .A(\EXU/_0558_ ), .B(\EXU/_0742_ ), .S(\EXU/_1082_ ), .Z(\EXU/_0243_ ) );
MUX2_X1 \EXU/_2237_ ( .A(\EXU/_0528_ ), .B(\EXU/_0712_ ), .S(\EXU/_1082_ ), .Z(\EXU/_0244_ ) );
MUX2_X1 \EXU/_2238_ ( .A(\EXU/_0529_ ), .B(\EXU/_0713_ ), .S(\EXU/_1082_ ), .Z(\EXU/_0245_ ) );
MUX2_X1 \EXU/_2239_ ( .A(\EXU/_0530_ ), .B(\EXU/_0714_ ), .S(\EXU/_1082_ ), .Z(\EXU/_0246_ ) );
MUX2_X1 \EXU/_2240_ ( .A(\EXU/_0531_ ), .B(\EXU/_0715_ ), .S(\EXU/_1082_ ), .Z(\EXU/_0247_ ) );
MUX2_X1 \EXU/_2241_ ( .A(\EXU/_0532_ ), .B(\EXU/_0716_ ), .S(\EXU/_1082_ ), .Z(\EXU/_0248_ ) );
BUF_X4 \EXU/_2242_ ( .A(\EXU/_1074_ ), .Z(\EXU/_1083_ ) );
MUX2_X1 \EXU/_2243_ ( .A(\EXU/_0533_ ), .B(\EXU/_0717_ ), .S(\EXU/_1083_ ), .Z(\EXU/_0249_ ) );
MUX2_X1 \EXU/_2244_ ( .A(\EXU/_0534_ ), .B(\EXU/_0718_ ), .S(\EXU/_1083_ ), .Z(\EXU/_0250_ ) );
MUX2_X1 \EXU/_2245_ ( .A(\EXU/_0535_ ), .B(\EXU/_0719_ ), .S(\EXU/_1083_ ), .Z(\EXU/_0251_ ) );
MUX2_X1 \EXU/_2246_ ( .A(\EXU/_0536_ ), .B(\EXU/_0720_ ), .S(\EXU/_1083_ ), .Z(\EXU/_0252_ ) );
MUX2_X1 \EXU/_2247_ ( .A(\EXU/_0537_ ), .B(\EXU/_0721_ ), .S(\EXU/_1083_ ), .Z(\EXU/_0253_ ) );
MUX2_X1 \EXU/_2248_ ( .A(\EXU/_0539_ ), .B(\EXU/_0723_ ), .S(\EXU/_1083_ ), .Z(\EXU/_0254_ ) );
MUX2_X1 \EXU/_2249_ ( .A(\EXU/_0540_ ), .B(\EXU/_0724_ ), .S(\EXU/_1083_ ), .Z(\EXU/_0255_ ) );
MUX2_X1 \EXU/_2250_ ( .A(\EXU/_0541_ ), .B(\EXU/_0725_ ), .S(\EXU/_1083_ ), .Z(\EXU/_0256_ ) );
MUX2_X1 \EXU/_2251_ ( .A(\EXU/_0542_ ), .B(\EXU/_0726_ ), .S(\EXU/_1083_ ), .Z(\EXU/_0257_ ) );
MUX2_X1 \EXU/_2252_ ( .A(\EXU/_0543_ ), .B(\EXU/_0727_ ), .S(\EXU/_1083_ ), .Z(\EXU/_0258_ ) );
BUF_X4 \EXU/_2253_ ( .A(\EXU/_1074_ ), .Z(\EXU/_1084_ ) );
MUX2_X1 \EXU/_2254_ ( .A(\EXU/_0544_ ), .B(\EXU/_0728_ ), .S(\EXU/_1084_ ), .Z(\EXU/_0259_ ) );
MUX2_X1 \EXU/_2255_ ( .A(\EXU/_0545_ ), .B(\EXU/_0729_ ), .S(\EXU/_1084_ ), .Z(\EXU/_0260_ ) );
MUX2_X1 \EXU/_2256_ ( .A(\EXU/_0546_ ), .B(\EXU/_0730_ ), .S(\EXU/_1084_ ), .Z(\EXU/_0261_ ) );
MUX2_X1 \EXU/_2257_ ( .A(\EXU/_0547_ ), .B(\EXU/_0731_ ), .S(\EXU/_1084_ ), .Z(\EXU/_0262_ ) );
MUX2_X1 \EXU/_2258_ ( .A(\EXU/_0548_ ), .B(\EXU/_0732_ ), .S(\EXU/_1084_ ), .Z(\EXU/_0263_ ) );
MUX2_X1 \EXU/_2259_ ( .A(\EXU/_0550_ ), .B(\EXU/_0734_ ), .S(\EXU/_1084_ ), .Z(\EXU/_0264_ ) );
MUX2_X1 \EXU/_2260_ ( .A(\EXU/_0551_ ), .B(\EXU/_0735_ ), .S(\EXU/_1084_ ), .Z(\EXU/_0265_ ) );
MUX2_X1 \EXU/_2261_ ( .A(\EXU/_0395_ ), .B(\EXU/_0615_ ), .S(\EXU/_1084_ ), .Z(\EXU/_0266_ ) );
MUX2_X1 \EXU/_2262_ ( .A(\EXU/_0406_ ), .B(\EXU/_0626_ ), .S(\EXU/_1084_ ), .Z(\EXU/_0267_ ) );
MUX2_X1 \EXU/_2263_ ( .A(\EXU/_0417_ ), .B(\EXU/_0637_ ), .S(\EXU/_1084_ ), .Z(\EXU/_0268_ ) );
BUF_X4 \EXU/_2264_ ( .A(\EXU/_1073_ ), .Z(\EXU/_1085_ ) );
MUX2_X1 \EXU/_2265_ ( .A(\EXU/_0420_ ), .B(\EXU/_0640_ ), .S(\EXU/_1085_ ), .Z(\EXU/_0269_ ) );
MUX2_X1 \EXU/_2266_ ( .A(\EXU/_0421_ ), .B(\EXU/_0641_ ), .S(\EXU/_1085_ ), .Z(\EXU/_0270_ ) );
MUX2_X1 \EXU/_2267_ ( .A(\EXU/_0422_ ), .B(\EXU/_0642_ ), .S(\EXU/_1085_ ), .Z(\EXU/_0271_ ) );
MUX2_X1 \EXU/_2268_ ( .A(\EXU/_0423_ ), .B(\EXU/_0643_ ), .S(\EXU/_1085_ ), .Z(\EXU/_0272_ ) );
MUX2_X1 \EXU/_2269_ ( .A(\EXU/_0424_ ), .B(\EXU/_0644_ ), .S(\EXU/_1085_ ), .Z(\EXU/_0273_ ) );
MUX2_X1 \EXU/_2270_ ( .A(\EXU/_0425_ ), .B(\EXU/_0645_ ), .S(\EXU/_1085_ ), .Z(\EXU/_0274_ ) );
MUX2_X1 \EXU/_2271_ ( .A(\EXU/_0426_ ), .B(\EXU/_0646_ ), .S(\EXU/_1085_ ), .Z(\EXU/_0275_ ) );
MUX2_X1 \EXU/_2272_ ( .A(\EXU/_0396_ ), .B(\EXU/_0616_ ), .S(\EXU/_1085_ ), .Z(\EXU/_0276_ ) );
MUX2_X1 \EXU/_2273_ ( .A(\EXU/_0397_ ), .B(\EXU/_0617_ ), .S(\EXU/_1085_ ), .Z(\EXU/_0277_ ) );
MUX2_X1 \EXU/_2274_ ( .A(\EXU/_0398_ ), .B(\EXU/_0618_ ), .S(\EXU/_1085_ ), .Z(\EXU/_0278_ ) );
BUF_X4 \EXU/_2275_ ( .A(\EXU/_1073_ ), .Z(\EXU/_1086_ ) );
MUX2_X1 \EXU/_2276_ ( .A(\EXU/_0399_ ), .B(\EXU/_0619_ ), .S(\EXU/_1086_ ), .Z(\EXU/_0279_ ) );
MUX2_X1 \EXU/_2277_ ( .A(\EXU/_0400_ ), .B(\EXU/_0620_ ), .S(\EXU/_1086_ ), .Z(\EXU/_0280_ ) );
MUX2_X1 \EXU/_2278_ ( .A(\EXU/_0401_ ), .B(\EXU/_0621_ ), .S(\EXU/_1086_ ), .Z(\EXU/_0281_ ) );
MUX2_X1 \EXU/_2279_ ( .A(\EXU/_0402_ ), .B(\EXU/_0622_ ), .S(\EXU/_1086_ ), .Z(\EXU/_0282_ ) );
MUX2_X1 \EXU/_2280_ ( .A(\EXU/_0403_ ), .B(\EXU/_0623_ ), .S(\EXU/_1086_ ), .Z(\EXU/_0283_ ) );
MUX2_X1 \EXU/_2281_ ( .A(\EXU/_0404_ ), .B(\EXU/_0624_ ), .S(\EXU/_1086_ ), .Z(\EXU/_0284_ ) );
MUX2_X1 \EXU/_2282_ ( .A(\EXU/_0405_ ), .B(\EXU/_0625_ ), .S(\EXU/_1086_ ), .Z(\EXU/_0285_ ) );
MUX2_X1 \EXU/_2283_ ( .A(\EXU/_0407_ ), .B(\EXU/_0627_ ), .S(\EXU/_1086_ ), .Z(\EXU/_0286_ ) );
MUX2_X1 \EXU/_2284_ ( .A(\EXU/_0408_ ), .B(\EXU/_0628_ ), .S(\EXU/_1086_ ), .Z(\EXU/_0287_ ) );
MUX2_X1 \EXU/_2285_ ( .A(\EXU/_0409_ ), .B(\EXU/_0629_ ), .S(\EXU/_1086_ ), .Z(\EXU/_0288_ ) );
BUF_X4 \EXU/_2286_ ( .A(\EXU/_1073_ ), .Z(\EXU/_1087_ ) );
MUX2_X1 \EXU/_2287_ ( .A(\EXU/_0410_ ), .B(\EXU/_0630_ ), .S(\EXU/_1087_ ), .Z(\EXU/_0289_ ) );
MUX2_X1 \EXU/_2288_ ( .A(\EXU/_0411_ ), .B(\EXU/_0631_ ), .S(\EXU/_1087_ ), .Z(\EXU/_0290_ ) );
MUX2_X1 \EXU/_2289_ ( .A(\EXU/_0412_ ), .B(\EXU/_0632_ ), .S(\EXU/_1087_ ), .Z(\EXU/_0291_ ) );
MUX2_X1 \EXU/_2290_ ( .A(\EXU/_0413_ ), .B(\EXU/_0633_ ), .S(\EXU/_1087_ ), .Z(\EXU/_0292_ ) );
MUX2_X1 \EXU/_2291_ ( .A(\EXU/_0414_ ), .B(\EXU/_0634_ ), .S(\EXU/_1087_ ), .Z(\EXU/_0293_ ) );
MUX2_X1 \EXU/_2292_ ( .A(\EXU/_0415_ ), .B(\EXU/_0635_ ), .S(\EXU/_1087_ ), .Z(\EXU/_0294_ ) );
MUX2_X1 \EXU/_2293_ ( .A(\EXU/_0416_ ), .B(\EXU/_0636_ ), .S(\EXU/_1087_ ), .Z(\EXU/_0295_ ) );
MUX2_X1 \EXU/_2294_ ( .A(\EXU/_0418_ ), .B(\EXU/_0638_ ), .S(\EXU/_1087_ ), .Z(\EXU/_0296_ ) );
MUX2_X1 \EXU/_2295_ ( .A(\EXU/_0419_ ), .B(\EXU/_0639_ ), .S(\EXU/_1087_ ), .Z(\EXU/_0297_ ) );
MUX2_X1 \EXU/_2296_ ( .A(\EXU/_0491_ ), .B(\EXU/_0743_ ), .S(\EXU/_1087_ ), .Z(\EXU/_0298_ ) );
BUF_X4 \EXU/_2297_ ( .A(\EXU/_1073_ ), .Z(\EXU/_1088_ ) );
MUX2_X1 \EXU/_2298_ ( .A(\EXU/_0502_ ), .B(\EXU/_0754_ ), .S(\EXU/_1088_ ), .Z(\EXU/_0299_ ) );
MUX2_X1 \EXU/_2299_ ( .A(\EXU/_0513_ ), .B(\EXU/_0765_ ), .S(\EXU/_1088_ ), .Z(\EXU/_0300_ ) );
MUX2_X1 \EXU/_2300_ ( .A(\EXU/_0516_ ), .B(\EXU/_0768_ ), .S(\EXU/_1088_ ), .Z(\EXU/_0301_ ) );
MUX2_X1 \EXU/_2301_ ( .A(\EXU/_0517_ ), .B(\EXU/_0769_ ), .S(\EXU/_1088_ ), .Z(\EXU/_0302_ ) );
MUX2_X1 \EXU/_2302_ ( .A(\EXU/_0518_ ), .B(\EXU/_0770_ ), .S(\EXU/_1088_ ), .Z(\EXU/_0303_ ) );
MUX2_X1 \EXU/_2303_ ( .A(\EXU/_0519_ ), .B(\EXU/_0771_ ), .S(\EXU/_1088_ ), .Z(\EXU/_0304_ ) );
MUX2_X1 \EXU/_2304_ ( .A(\EXU/_0520_ ), .B(\EXU/_0772_ ), .S(\EXU/_1088_ ), .Z(\EXU/_0305_ ) );
MUX2_X1 \EXU/_2305_ ( .A(\EXU/_0521_ ), .B(\EXU/_0773_ ), .S(\EXU/_1088_ ), .Z(\EXU/_0306_ ) );
MUX2_X1 \EXU/_2306_ ( .A(\EXU/_0522_ ), .B(\EXU/_0774_ ), .S(\EXU/_1088_ ), .Z(\EXU/_0307_ ) );
MUX2_X1 \EXU/_2307_ ( .A(\EXU/_0492_ ), .B(\EXU/_0744_ ), .S(\EXU/_1088_ ), .Z(\EXU/_0308_ ) );
BUF_X4 \EXU/_2308_ ( .A(\EXU/_1073_ ), .Z(\EXU/_1089_ ) );
MUX2_X1 \EXU/_2309_ ( .A(\EXU/_0493_ ), .B(\EXU/_0745_ ), .S(\EXU/_1089_ ), .Z(\EXU/_0309_ ) );
MUX2_X1 \EXU/_2310_ ( .A(\EXU/_0494_ ), .B(\EXU/_0746_ ), .S(\EXU/_1089_ ), .Z(\EXU/_0310_ ) );
MUX2_X1 \EXU/_2311_ ( .A(\EXU/_0495_ ), .B(\EXU/_0747_ ), .S(\EXU/_1089_ ), .Z(\EXU/_0311_ ) );
MUX2_X1 \EXU/_2312_ ( .A(\EXU/_0496_ ), .B(\EXU/_0748_ ), .S(\EXU/_1089_ ), .Z(\EXU/_0312_ ) );
MUX2_X1 \EXU/_2313_ ( .A(\EXU/_0497_ ), .B(\EXU/_0749_ ), .S(\EXU/_1089_ ), .Z(\EXU/_0313_ ) );
MUX2_X1 \EXU/_2314_ ( .A(\EXU/_0498_ ), .B(\EXU/_0750_ ), .S(\EXU/_1089_ ), .Z(\EXU/_0314_ ) );
MUX2_X1 \EXU/_2315_ ( .A(\EXU/_0499_ ), .B(\EXU/_0751_ ), .S(\EXU/_1089_ ), .Z(\EXU/_0315_ ) );
MUX2_X1 \EXU/_2316_ ( .A(\EXU/_0500_ ), .B(\EXU/_0752_ ), .S(\EXU/_1089_ ), .Z(\EXU/_0316_ ) );
MUX2_X1 \EXU/_2317_ ( .A(\EXU/_0501_ ), .B(\EXU/_0753_ ), .S(\EXU/_1089_ ), .Z(\EXU/_0317_ ) );
MUX2_X1 \EXU/_2318_ ( .A(\EXU/_0503_ ), .B(\EXU/_0755_ ), .S(\EXU/_1089_ ), .Z(\EXU/_0318_ ) );
BUF_X4 \EXU/_2319_ ( .A(\EXU/_1073_ ), .Z(\EXU/_1090_ ) );
MUX2_X1 \EXU/_2320_ ( .A(\EXU/_0504_ ), .B(\EXU/_0756_ ), .S(\EXU/_1090_ ), .Z(\EXU/_0319_ ) );
MUX2_X1 \EXU/_2321_ ( .A(\EXU/_0505_ ), .B(\EXU/_0757_ ), .S(\EXU/_1090_ ), .Z(\EXU/_0320_ ) );
MUX2_X1 \EXU/_2322_ ( .A(\EXU/_0506_ ), .B(\EXU/_0758_ ), .S(\EXU/_1090_ ), .Z(\EXU/_0321_ ) );
MUX2_X1 \EXU/_2323_ ( .A(\EXU/_0507_ ), .B(\EXU/_0759_ ), .S(\EXU/_1090_ ), .Z(\EXU/_0322_ ) );
MUX2_X1 \EXU/_2324_ ( .A(\EXU/_0508_ ), .B(\EXU/_0760_ ), .S(\EXU/_1090_ ), .Z(\EXU/_0323_ ) );
MUX2_X1 \EXU/_2325_ ( .A(\EXU/_0509_ ), .B(\EXU/_0761_ ), .S(\EXU/_1090_ ), .Z(\EXU/_0324_ ) );
MUX2_X1 \EXU/_2326_ ( .A(\EXU/_0510_ ), .B(\EXU/_0762_ ), .S(\EXU/_1090_ ), .Z(\EXU/_0325_ ) );
MUX2_X1 \EXU/_2327_ ( .A(\EXU/_0511_ ), .B(\EXU/_0763_ ), .S(\EXU/_1090_ ), .Z(\EXU/_0326_ ) );
MUX2_X1 \EXU/_2328_ ( .A(\EXU/_0512_ ), .B(\EXU/_0764_ ), .S(\EXU/_1090_ ), .Z(\EXU/_0327_ ) );
MUX2_X1 \EXU/_2329_ ( .A(\EXU/_0514_ ), .B(\EXU/_0766_ ), .S(\EXU/_1090_ ), .Z(\EXU/_0328_ ) );
BUF_X4 \EXU/_2330_ ( .A(\EXU/_1073_ ), .Z(\EXU/_1091_ ) );
MUX2_X1 \EXU/_2331_ ( .A(\EXU/_0515_ ), .B(\EXU/_0767_ ), .S(\EXU/_1091_ ), .Z(\EXU/_0329_ ) );
MUX2_X1 \EXU/_2332_ ( .A(\EXU/_0381_ ), .B(\EXU/_0596_ ), .S(\EXU/_1091_ ), .Z(\EXU/_0330_ ) );
MUX2_X1 \EXU/_2333_ ( .A(\EXU/_0382_ ), .B(\EXU/_0597_ ), .S(\EXU/_1091_ ), .Z(\EXU/_0331_ ) );
MUX2_X1 \EXU/_2334_ ( .A(\EXU/_0383_ ), .B(\EXU/_0598_ ), .S(\EXU/_1091_ ), .Z(\EXU/_0332_ ) );
MUX2_X1 \EXU/_2335_ ( .A(\EXU/_0384_ ), .B(\EXU/_0599_ ), .S(\EXU/_1091_ ), .Z(\EXU/_0333_ ) );
MUX2_X1 \EXU/_2336_ ( .A(\EXU/_0385_ ), .B(\EXU/_0600_ ), .S(\EXU/_1091_ ), .Z(\EXU/_0334_ ) );
MUX2_X1 \EXU/_2337_ ( .A(\EXU/_0386_ ), .B(\EXU/_0601_ ), .S(\EXU/_1091_ ), .Z(\EXU/_0335_ ) );
MUX2_X1 \EXU/_2338_ ( .A(\EXU/_0387_ ), .B(\EXU/_0602_ ), .S(\EXU/_1091_ ), .Z(\EXU/_0336_ ) );
MUX2_X1 \EXU/_2339_ ( .A(\EXU/_0394_ ), .B(\EXU/_0609_ ), .S(\EXU/_1091_ ), .Z(\EXU/_0337_ ) );
MUX2_X1 \EXU/_2340_ ( .A(\EXU/_0391_ ), .B(\EXU/_0606_ ), .S(\EXU/_1091_ ), .Z(\EXU/_0338_ ) );
BUF_X4 \EXU/_2341_ ( .A(\EXU/_1073_ ), .Z(\EXU/_1092_ ) );
MUX2_X1 \EXU/_2342_ ( .A(\EXU/_0392_ ), .B(\EXU/_0607_ ), .S(\EXU/_1092_ ), .Z(\EXU/_0339_ ) );
MUX2_X1 \EXU/_2343_ ( .A(\EXU/_0393_ ), .B(\EXU/_0608_ ), .S(\EXU/_1092_ ), .Z(\EXU/_0340_ ) );
MUX2_X1 \EXU/_2344_ ( .A(\EXU/_0388_ ), .B(\EXU/_0603_ ), .S(\EXU/_1092_ ), .Z(\EXU/_0341_ ) );
MUX2_X1 \EXU/_2345_ ( .A(\EXU/_0389_ ), .B(\EXU/_0604_ ), .S(\EXU/_1092_ ), .Z(\EXU/_0342_ ) );
MUX2_X1 \EXU/_2346_ ( .A(\EXU/_0390_ ), .B(\EXU/_0605_ ), .S(\EXU/_1092_ ), .Z(\EXU/_0343_ ) );
MUX2_X1 \EXU/_2347_ ( .A(\EXU/_0526_ ), .B(\EXU/_0613_ ), .S(\EXU/_1092_ ), .Z(\EXU/_0344_ ) );
MUX2_X1 \EXU/_2348_ ( .A(\EXU/_0559_ ), .B(\EXU/_0614_ ), .S(\EXU/_1092_ ), .Z(\EXU/_0345_ ) );
MUX2_X1 \EXU/_2349_ ( .A(\EXU/_0523_ ), .B(\EXU/_0610_ ), .S(\EXU/_1092_ ), .Z(\EXU/_0346_ ) );
MUX2_X1 \EXU/_2350_ ( .A(\EXU/_0524_ ), .B(\EXU/_0611_ ), .S(\EXU/_1092_ ), .Z(\EXU/_0347_ ) );
MUX2_X1 \EXU/_2351_ ( .A(\EXU/_0525_ ), .B(\EXU/_0612_ ), .S(\EXU/_1092_ ), .Z(\EXU/_0348_ ) );
NOR3_X1 \EXU/_2352_ ( .A1(\EXU/_1101_ ), .A2(\EXU/_1216_ ), .A3(\EXU/_0560_ ), .ZN(\EXU/_1093_ ) );
NOR3_X1 \EXU/_2353_ ( .A1(\EXU/_1069_ ), .A2(\EXU/_1075_ ), .A3(\EXU/_1093_ ), .ZN(\EXU/_1094_ ) );
NAND3_X1 \EXU/_2354_ ( .A1(\EXU/_1215_ ), .A2(\EXU/_1216_ ), .A3(\EXU/_0841_ ), .ZN(\EXU/_1095_ ) );
AND2_X1 \EXU/_2355_ ( .A1(\EXU/_0842_ ), .A2(\EXU/_1095_ ), .ZN(\EXU/_1096_ ) );
INV_X1 \EXU/_2356_ ( .A(\EXU/_1096_ ), .ZN(\EXU/_1097_ ) );
AOI21_X1 \EXU/_2357_ ( .A(\EXU/_1214_ ), .B1(\EXU/_1094_ ), .B2(\EXU/_1097_ ), .ZN(\EXU/_0168_ ) );
INV_X1 \EXU/_2358_ ( .A(\EXU/_1073_ ), .ZN(\EXU/_1098_ ) );
NOR3_X1 \EXU/_2359_ ( .A1(\EXU/_1098_ ), .A2(\EXU/_0613_ ), .A3(\EXU/_0614_ ), .ZN(\EXU/_1099_ ) );
AOI211_X4 \EXU/_2360_ ( .A(\EXU/_0594_ ), .B(\EXU/_1099_ ), .C1(\EXU/_0560_ ), .C2(\EXU/_0561_ ), .ZN(\EXU/_1100_ ) );
AOI21_X1 \EXU/_2361_ ( .A(\EXU/_1214_ ), .B1(\EXU/_1100_ ), .B2(\EXU/_1097_ ), .ZN(\EXU/_0169_ ) );
DFF_X1 \EXU/_2362_ ( .D(\EXU/_1430_ ), .CK(clock ), .Q(\_EXU_io_out_bits_memOut [0] ), .QN(\EXU/_1429_ ) );
DFF_X1 \EXU/_2363_ ( .D(\EXU/_1431_ ), .CK(clock ), .Q(\_EXU_io_out_bits_memOut [1] ), .QN(\EXU/_1428_ ) );
DFF_X1 \EXU/_2364_ ( .D(\EXU/_1432_ ), .CK(clock ), .Q(\_EXU_io_out_bits_memOut [2] ), .QN(\EXU/_1427_ ) );
DFF_X1 \EXU/_2365_ ( .D(\EXU/_1433_ ), .CK(clock ), .Q(\_EXU_io_out_bits_memOut [3] ), .QN(\EXU/_1426_ ) );
DFF_X1 \EXU/_2366_ ( .D(\EXU/_1434_ ), .CK(clock ), .Q(\_EXU_io_out_bits_memOut [4] ), .QN(\EXU/_1425_ ) );
DFF_X1 \EXU/_2367_ ( .D(\EXU/_1435_ ), .CK(clock ), .Q(\_EXU_io_out_bits_memOut [5] ), .QN(\EXU/_1424_ ) );
DFF_X1 \EXU/_2368_ ( .D(\EXU/_1436_ ), .CK(clock ), .Q(\_EXU_io_out_bits_memOut [6] ), .QN(\EXU/_1423_ ) );
DFF_X1 \EXU/_2369_ ( .D(\EXU/_1437_ ), .CK(clock ), .Q(\_EXU_io_out_bits_memOut [7] ), .QN(\EXU/_1422_ ) );
DFF_X1 \EXU/_2370_ ( .D(\EXU/_1438_ ), .CK(clock ), .Q(\_EXU_io_out_bits_memOut [8] ), .QN(\EXU/_1421_ ) );
DFF_X1 \EXU/_2371_ ( .D(\EXU/_1439_ ), .CK(clock ), .Q(\_EXU_io_out_bits_memOut [9] ), .QN(\EXU/_1420_ ) );
DFF_X1 \EXU/_2372_ ( .D(\EXU/_1440_ ), .CK(clock ), .Q(\_EXU_io_out_bits_memOut [10] ), .QN(\EXU/_1419_ ) );
DFF_X1 \EXU/_2373_ ( .D(\EXU/_1441_ ), .CK(clock ), .Q(\_EXU_io_out_bits_memOut [11] ), .QN(\EXU/_1418_ ) );
DFF_X1 \EXU/_2374_ ( .D(\EXU/_1442_ ), .CK(clock ), .Q(\_EXU_io_out_bits_memOut [12] ), .QN(\EXU/_1417_ ) );
DFF_X1 \EXU/_2375_ ( .D(\EXU/_1443_ ), .CK(clock ), .Q(\_EXU_io_out_bits_memOut [13] ), .QN(\EXU/_1416_ ) );
DFF_X1 \EXU/_2376_ ( .D(\EXU/_1444_ ), .CK(clock ), .Q(\_EXU_io_out_bits_memOut [14] ), .QN(\EXU/_1415_ ) );
DFF_X1 \EXU/_2377_ ( .D(\EXU/_1445_ ), .CK(clock ), .Q(\_EXU_io_out_bits_memOut [15] ), .QN(\EXU/_1414_ ) );
DFF_X1 \EXU/_2378_ ( .D(\EXU/_1446_ ), .CK(clock ), .Q(\_EXU_io_out_bits_memOut [16] ), .QN(\EXU/_1413_ ) );
DFF_X1 \EXU/_2379_ ( .D(\EXU/_1447_ ), .CK(clock ), .Q(\_EXU_io_out_bits_memOut [17] ), .QN(\EXU/_1412_ ) );
DFF_X1 \EXU/_2380_ ( .D(\EXU/_1448_ ), .CK(clock ), .Q(\_EXU_io_out_bits_memOut [18] ), .QN(\EXU/_1411_ ) );
DFF_X1 \EXU/_2381_ ( .D(\EXU/_1449_ ), .CK(clock ), .Q(\_EXU_io_out_bits_memOut [19] ), .QN(\EXU/_1410_ ) );
DFF_X1 \EXU/_2382_ ( .D(\EXU/_1450_ ), .CK(clock ), .Q(\_EXU_io_out_bits_memOut [20] ), .QN(\EXU/_1409_ ) );
DFF_X1 \EXU/_2383_ ( .D(\EXU/_1451_ ), .CK(clock ), .Q(\_EXU_io_out_bits_memOut [21] ), .QN(\EXU/_1408_ ) );
DFF_X1 \EXU/_2384_ ( .D(\EXU/_1452_ ), .CK(clock ), .Q(\_EXU_io_out_bits_memOut [22] ), .QN(\EXU/_1407_ ) );
DFF_X1 \EXU/_2385_ ( .D(\EXU/_1453_ ), .CK(clock ), .Q(\_EXU_io_out_bits_memOut [23] ), .QN(\EXU/_1406_ ) );
DFF_X1 \EXU/_2386_ ( .D(\EXU/_1454_ ), .CK(clock ), .Q(\_EXU_io_out_bits_memOut [24] ), .QN(\EXU/_1405_ ) );
DFF_X1 \EXU/_2387_ ( .D(\EXU/_1455_ ), .CK(clock ), .Q(\_EXU_io_out_bits_memOut [25] ), .QN(\EXU/_1404_ ) );
DFF_X1 \EXU/_2388_ ( .D(\EXU/_1456_ ), .CK(clock ), .Q(\_EXU_io_out_bits_memOut [26] ), .QN(\EXU/_1403_ ) );
DFF_X1 \EXU/_2389_ ( .D(\EXU/_1457_ ), .CK(clock ), .Q(\_EXU_io_out_bits_memOut [27] ), .QN(\EXU/_1402_ ) );
DFF_X1 \EXU/_2390_ ( .D(\EXU/_1458_ ), .CK(clock ), .Q(\_EXU_io_out_bits_memOut [28] ), .QN(\EXU/_1401_ ) );
DFF_X1 \EXU/_2391_ ( .D(\EXU/_1459_ ), .CK(clock ), .Q(\_EXU_io_out_bits_memOut [29] ), .QN(\EXU/_1400_ ) );
DFF_X1 \EXU/_2392_ ( .D(\EXU/_1460_ ), .CK(clock ), .Q(\_EXU_io_out_bits_memOut [30] ), .QN(\EXU/_1399_ ) );
DFF_X1 \EXU/_2393_ ( .D(\EXU/_1461_ ), .CK(clock ), .Q(\_EXU_io_out_bits_memOut [31] ), .QN(\EXU/_1398_ ) );
DFF_X1 \EXU/_2394_ ( .D(\EXU/_1462_ ), .CK(clock ), .Q(\EXU/state [0] ), .QN(\EXU/_1397_ ) );
DFF_X1 \EXU/_2395_ ( .D(\EXU/_1463_ ), .CK(clock ), .Q(\EXU/state [1] ), .QN(\EXU/_1396_ ) );
DFF_X1 \EXU/_2396_ ( .D(\EXU/_1464_ ), .CK(clock ), .Q(\EXU/in_pc [0] ), .QN(\EXU/_1395_ ) );
DFF_X1 \EXU/_2397_ ( .D(\EXU/_1465_ ), .CK(clock ), .Q(\EXU/in_pc [1] ), .QN(\EXU/_1394_ ) );
DFF_X1 \EXU/_2398_ ( .D(\EXU/_1466_ ), .CK(clock ), .Q(\EXU/in_pc [2] ), .QN(\EXU/_1393_ ) );
DFF_X1 \EXU/_2399_ ( .D(\EXU/_1467_ ), .CK(clock ), .Q(\EXU/in_pc [3] ), .QN(\EXU/_1392_ ) );
DFF_X1 \EXU/_2400_ ( .D(\EXU/_1468_ ), .CK(clock ), .Q(\EXU/in_pc [4] ), .QN(\EXU/_1391_ ) );
DFF_X1 \EXU/_2401_ ( .D(\EXU/_1469_ ), .CK(clock ), .Q(\EXU/in_pc [5] ), .QN(\EXU/_1390_ ) );
DFF_X1 \EXU/_2402_ ( .D(\EXU/_1470_ ), .CK(clock ), .Q(\EXU/in_pc [6] ), .QN(\EXU/_1389_ ) );
DFF_X1 \EXU/_2403_ ( .D(\EXU/_1471_ ), .CK(clock ), .Q(\EXU/in_pc [7] ), .QN(\EXU/_1388_ ) );
DFF_X1 \EXU/_2404_ ( .D(\EXU/_1472_ ), .CK(clock ), .Q(\EXU/in_pc [8] ), .QN(\EXU/_1387_ ) );
DFF_X1 \EXU/_2405_ ( .D(\EXU/_1473_ ), .CK(clock ), .Q(\EXU/in_pc [9] ), .QN(\EXU/_1386_ ) );
DFF_X1 \EXU/_2406_ ( .D(\EXU/_1474_ ), .CK(clock ), .Q(\EXU/in_pc [10] ), .QN(\EXU/_1385_ ) );
DFF_X1 \EXU/_2407_ ( .D(\EXU/_1475_ ), .CK(clock ), .Q(\EXU/in_pc [11] ), .QN(\EXU/_1384_ ) );
DFF_X1 \EXU/_2408_ ( .D(\EXU/_1476_ ), .CK(clock ), .Q(\EXU/in_pc [12] ), .QN(\EXU/_1383_ ) );
DFF_X1 \EXU/_2409_ ( .D(\EXU/_1477_ ), .CK(clock ), .Q(\EXU/in_pc [13] ), .QN(\EXU/_1382_ ) );
DFF_X1 \EXU/_2410_ ( .D(\EXU/_1478_ ), .CK(clock ), .Q(\EXU/in_pc [14] ), .QN(\EXU/_1381_ ) );
DFF_X1 \EXU/_2411_ ( .D(\EXU/_1479_ ), .CK(clock ), .Q(\EXU/in_pc [15] ), .QN(\EXU/_1380_ ) );
DFF_X1 \EXU/_2412_ ( .D(\EXU/_1480_ ), .CK(clock ), .Q(\EXU/in_pc [16] ), .QN(\EXU/_1379_ ) );
DFF_X1 \EXU/_2413_ ( .D(\EXU/_1481_ ), .CK(clock ), .Q(\EXU/in_pc [17] ), .QN(\EXU/_1378_ ) );
DFF_X1 \EXU/_2414_ ( .D(\EXU/_1482_ ), .CK(clock ), .Q(\EXU/in_pc [18] ), .QN(\EXU/_1377_ ) );
DFF_X1 \EXU/_2415_ ( .D(\EXU/_1483_ ), .CK(clock ), .Q(\EXU/in_pc [19] ), .QN(\EXU/_1376_ ) );
DFF_X1 \EXU/_2416_ ( .D(\EXU/_1484_ ), .CK(clock ), .Q(\EXU/in_pc [20] ), .QN(\EXU/_1375_ ) );
DFF_X1 \EXU/_2417_ ( .D(\EXU/_1485_ ), .CK(clock ), .Q(\EXU/in_pc [21] ), .QN(\EXU/_1374_ ) );
DFF_X1 \EXU/_2418_ ( .D(\EXU/_1486_ ), .CK(clock ), .Q(\EXU/in_pc [22] ), .QN(\EXU/_1373_ ) );
DFF_X1 \EXU/_2419_ ( .D(\EXU/_1487_ ), .CK(clock ), .Q(\EXU/in_pc [23] ), .QN(\EXU/_1372_ ) );
DFF_X1 \EXU/_2420_ ( .D(\EXU/_1488_ ), .CK(clock ), .Q(\EXU/in_pc [24] ), .QN(\EXU/_1371_ ) );
DFF_X1 \EXU/_2421_ ( .D(\EXU/_1489_ ), .CK(clock ), .Q(\EXU/in_pc [25] ), .QN(\EXU/_1370_ ) );
DFF_X1 \EXU/_2422_ ( .D(\EXU/_1490_ ), .CK(clock ), .Q(\EXU/in_pc [26] ), .QN(\EXU/_1369_ ) );
DFF_X1 \EXU/_2423_ ( .D(\EXU/_1491_ ), .CK(clock ), .Q(\EXU/in_pc [27] ), .QN(\EXU/_1368_ ) );
DFF_X1 \EXU/_2424_ ( .D(\EXU/_1492_ ), .CK(clock ), .Q(\EXU/in_pc [28] ), .QN(\EXU/_1367_ ) );
DFF_X1 \EXU/_2425_ ( .D(\EXU/_1493_ ), .CK(clock ), .Q(\EXU/in_pc [29] ), .QN(\EXU/_1366_ ) );
DFF_X1 \EXU/_2426_ ( .D(\EXU/_1494_ ), .CK(clock ), .Q(\EXU/in_pc [30] ), .QN(\EXU/_1365_ ) );
DFF_X1 \EXU/_2427_ ( .D(\EXU/_1495_ ), .CK(clock ), .Q(\EXU/in_pc [31] ), .QN(\EXU/_1364_ ) );
DFF_X1 \EXU/_2428_ ( .D(\EXU/_1496_ ), .CK(clock ), .Q(\EXU/in_rd1 [0] ), .QN(\EXU/_1363_ ) );
DFF_X1 \EXU/_2429_ ( .D(\EXU/_1497_ ), .CK(clock ), .Q(\EXU/in_rd1 [1] ), .QN(\EXU/_1362_ ) );
DFF_X1 \EXU/_2430_ ( .D(\EXU/_1498_ ), .CK(clock ), .Q(\EXU/in_rd1 [2] ), .QN(\EXU/_1361_ ) );
DFF_X1 \EXU/_2431_ ( .D(\EXU/_1499_ ), .CK(clock ), .Q(\EXU/in_rd1 [3] ), .QN(\EXU/_1360_ ) );
DFF_X1 \EXU/_2432_ ( .D(\EXU/_1500_ ), .CK(clock ), .Q(\EXU/in_rd1 [4] ), .QN(\EXU/_1359_ ) );
DFF_X1 \EXU/_2433_ ( .D(\EXU/_1501_ ), .CK(clock ), .Q(\EXU/in_rd1 [5] ), .QN(\EXU/_1358_ ) );
DFF_X1 \EXU/_2434_ ( .D(\EXU/_1502_ ), .CK(clock ), .Q(\EXU/in_rd1 [6] ), .QN(\EXU/_1357_ ) );
DFF_X1 \EXU/_2435_ ( .D(\EXU/_1503_ ), .CK(clock ), .Q(\EXU/in_rd1 [7] ), .QN(\EXU/_1356_ ) );
DFF_X1 \EXU/_2436_ ( .D(\EXU/_1504_ ), .CK(clock ), .Q(\EXU/in_rd1 [8] ), .QN(\EXU/_1355_ ) );
DFF_X1 \EXU/_2437_ ( .D(\EXU/_1505_ ), .CK(clock ), .Q(\EXU/in_rd1 [9] ), .QN(\EXU/_1354_ ) );
DFF_X1 \EXU/_2438_ ( .D(\EXU/_1506_ ), .CK(clock ), .Q(\EXU/in_rd1 [10] ), .QN(\EXU/_1353_ ) );
DFF_X1 \EXU/_2439_ ( .D(\EXU/_1507_ ), .CK(clock ), .Q(\EXU/in_rd1 [11] ), .QN(\EXU/_1352_ ) );
DFF_X1 \EXU/_2440_ ( .D(\EXU/_1508_ ), .CK(clock ), .Q(\EXU/in_rd1 [12] ), .QN(\EXU/_1351_ ) );
DFF_X1 \EXU/_2441_ ( .D(\EXU/_1509_ ), .CK(clock ), .Q(\EXU/in_rd1 [13] ), .QN(\EXU/_1350_ ) );
DFF_X1 \EXU/_2442_ ( .D(\EXU/_1510_ ), .CK(clock ), .Q(\EXU/in_rd1 [14] ), .QN(\EXU/_1349_ ) );
DFF_X1 \EXU/_2443_ ( .D(\EXU/_1511_ ), .CK(clock ), .Q(\EXU/in_rd1 [15] ), .QN(\EXU/_1348_ ) );
DFF_X1 \EXU/_2444_ ( .D(\EXU/_1512_ ), .CK(clock ), .Q(\EXU/in_rd1 [16] ), .QN(\EXU/_1347_ ) );
DFF_X1 \EXU/_2445_ ( .D(\EXU/_1513_ ), .CK(clock ), .Q(\EXU/in_rd1 [17] ), .QN(\EXU/_1346_ ) );
DFF_X1 \EXU/_2446_ ( .D(\EXU/_1514_ ), .CK(clock ), .Q(\EXU/in_rd1 [18] ), .QN(\EXU/_1345_ ) );
DFF_X1 \EXU/_2447_ ( .D(\EXU/_1515_ ), .CK(clock ), .Q(\EXU/in_rd1 [19] ), .QN(\EXU/_1344_ ) );
DFF_X1 \EXU/_2448_ ( .D(\EXU/_1516_ ), .CK(clock ), .Q(\EXU/in_rd1 [20] ), .QN(\EXU/_1343_ ) );
DFF_X1 \EXU/_2449_ ( .D(\EXU/_1517_ ), .CK(clock ), .Q(\EXU/in_rd1 [21] ), .QN(\EXU/_1342_ ) );
DFF_X1 \EXU/_2450_ ( .D(\EXU/_1518_ ), .CK(clock ), .Q(\EXU/in_rd1 [22] ), .QN(\EXU/_1341_ ) );
DFF_X1 \EXU/_2451_ ( .D(\EXU/_1519_ ), .CK(clock ), .Q(\EXU/in_rd1 [23] ), .QN(\EXU/_1340_ ) );
DFF_X1 \EXU/_2452_ ( .D(\EXU/_1520_ ), .CK(clock ), .Q(\EXU/in_rd1 [24] ), .QN(\EXU/_1339_ ) );
DFF_X1 \EXU/_2453_ ( .D(\EXU/_1521_ ), .CK(clock ), .Q(\EXU/in_rd1 [25] ), .QN(\EXU/_1338_ ) );
DFF_X1 \EXU/_2454_ ( .D(\EXU/_1522_ ), .CK(clock ), .Q(\EXU/in_rd1 [26] ), .QN(\EXU/_1337_ ) );
DFF_X1 \EXU/_2455_ ( .D(\EXU/_1523_ ), .CK(clock ), .Q(\EXU/in_rd1 [27] ), .QN(\EXU/_1336_ ) );
DFF_X1 \EXU/_2456_ ( .D(\EXU/_1524_ ), .CK(clock ), .Q(\EXU/in_rd1 [28] ), .QN(\EXU/_1335_ ) );
DFF_X1 \EXU/_2457_ ( .D(\EXU/_1525_ ), .CK(clock ), .Q(\EXU/in_rd1 [29] ), .QN(\EXU/_1334_ ) );
DFF_X1 \EXU/_2458_ ( .D(\EXU/_1526_ ), .CK(clock ), .Q(\EXU/in_rd1 [30] ), .QN(\EXU/_1333_ ) );
DFF_X1 \EXU/_2459_ ( .D(\EXU/_1527_ ), .CK(clock ), .Q(\EXU/in_rd1 [31] ), .QN(\EXU/_1332_ ) );
DFF_X1 \EXU/_2460_ ( .D(\EXU/_1528_ ), .CK(clock ), .Q(\_EXU_io_LSUIn_bits_wdata [0] ), .QN(\EXU/_1331_ ) );
DFF_X1 \EXU/_2461_ ( .D(\EXU/_1529_ ), .CK(clock ), .Q(\_EXU_io_LSUIn_bits_wdata [1] ), .QN(\EXU/_1330_ ) );
DFF_X1 \EXU/_2462_ ( .D(\EXU/_1530_ ), .CK(clock ), .Q(\_EXU_io_LSUIn_bits_wdata [2] ), .QN(\EXU/_1329_ ) );
DFF_X1 \EXU/_2463_ ( .D(\EXU/_1531_ ), .CK(clock ), .Q(\_EXU_io_LSUIn_bits_wdata [3] ), .QN(\EXU/_1328_ ) );
DFF_X1 \EXU/_2464_ ( .D(\EXU/_1532_ ), .CK(clock ), .Q(\_EXU_io_LSUIn_bits_wdata [4] ), .QN(\EXU/_1327_ ) );
DFF_X1 \EXU/_2465_ ( .D(\EXU/_1533_ ), .CK(clock ), .Q(\_EXU_io_LSUIn_bits_wdata [5] ), .QN(\EXU/_1326_ ) );
DFF_X1 \EXU/_2466_ ( .D(\EXU/_1534_ ), .CK(clock ), .Q(\_EXU_io_LSUIn_bits_wdata [6] ), .QN(\EXU/_1325_ ) );
DFF_X1 \EXU/_2467_ ( .D(\EXU/_1535_ ), .CK(clock ), .Q(\_EXU_io_LSUIn_bits_wdata [7] ), .QN(\EXU/_1324_ ) );
DFF_X1 \EXU/_2468_ ( .D(\EXU/_1536_ ), .CK(clock ), .Q(\_EXU_io_LSUIn_bits_wdata [8] ), .QN(\EXU/_1323_ ) );
DFF_X1 \EXU/_2469_ ( .D(\EXU/_1537_ ), .CK(clock ), .Q(\_EXU_io_LSUIn_bits_wdata [9] ), .QN(\EXU/_1322_ ) );
DFF_X1 \EXU/_2470_ ( .D(\EXU/_1538_ ), .CK(clock ), .Q(\_EXU_io_LSUIn_bits_wdata [10] ), .QN(\EXU/_1321_ ) );
DFF_X1 \EXU/_2471_ ( .D(\EXU/_1539_ ), .CK(clock ), .Q(\_EXU_io_LSUIn_bits_wdata [11] ), .QN(\EXU/_1320_ ) );
DFF_X1 \EXU/_2472_ ( .D(\EXU/_1540_ ), .CK(clock ), .Q(\_EXU_io_LSUIn_bits_wdata [12] ), .QN(\EXU/_1319_ ) );
DFF_X1 \EXU/_2473_ ( .D(\EXU/_1541_ ), .CK(clock ), .Q(\_EXU_io_LSUIn_bits_wdata [13] ), .QN(\EXU/_1318_ ) );
DFF_X1 \EXU/_2474_ ( .D(\EXU/_1542_ ), .CK(clock ), .Q(\_EXU_io_LSUIn_bits_wdata [14] ), .QN(\EXU/_1317_ ) );
DFF_X1 \EXU/_2475_ ( .D(\EXU/_1543_ ), .CK(clock ), .Q(\_EXU_io_LSUIn_bits_wdata [15] ), .QN(\EXU/_1316_ ) );
DFF_X1 \EXU/_2476_ ( .D(\EXU/_1544_ ), .CK(clock ), .Q(\_EXU_io_LSUIn_bits_wdata [16] ), .QN(\EXU/_1315_ ) );
DFF_X1 \EXU/_2477_ ( .D(\EXU/_1545_ ), .CK(clock ), .Q(\_EXU_io_LSUIn_bits_wdata [17] ), .QN(\EXU/_1314_ ) );
DFF_X1 \EXU/_2478_ ( .D(\EXU/_1546_ ), .CK(clock ), .Q(\_EXU_io_LSUIn_bits_wdata [18] ), .QN(\EXU/_1313_ ) );
DFF_X1 \EXU/_2479_ ( .D(\EXU/_1547_ ), .CK(clock ), .Q(\_EXU_io_LSUIn_bits_wdata [19] ), .QN(\EXU/_1312_ ) );
DFF_X1 \EXU/_2480_ ( .D(\EXU/_1548_ ), .CK(clock ), .Q(\_EXU_io_LSUIn_bits_wdata [20] ), .QN(\EXU/_1311_ ) );
DFF_X1 \EXU/_2481_ ( .D(\EXU/_1549_ ), .CK(clock ), .Q(\_EXU_io_LSUIn_bits_wdata [21] ), .QN(\EXU/_1310_ ) );
DFF_X1 \EXU/_2482_ ( .D(\EXU/_1550_ ), .CK(clock ), .Q(\_EXU_io_LSUIn_bits_wdata [22] ), .QN(\EXU/_1309_ ) );
DFF_X1 \EXU/_2483_ ( .D(\EXU/_1551_ ), .CK(clock ), .Q(\_EXU_io_LSUIn_bits_wdata [23] ), .QN(\EXU/_1308_ ) );
DFF_X1 \EXU/_2484_ ( .D(\EXU/_1552_ ), .CK(clock ), .Q(\_EXU_io_LSUIn_bits_wdata [24] ), .QN(\EXU/_1307_ ) );
DFF_X1 \EXU/_2485_ ( .D(\EXU/_1553_ ), .CK(clock ), .Q(\_EXU_io_LSUIn_bits_wdata [25] ), .QN(\EXU/_1306_ ) );
DFF_X1 \EXU/_2486_ ( .D(\EXU/_1554_ ), .CK(clock ), .Q(\_EXU_io_LSUIn_bits_wdata [26] ), .QN(\EXU/_1305_ ) );
DFF_X1 \EXU/_2487_ ( .D(\EXU/_1555_ ), .CK(clock ), .Q(\_EXU_io_LSUIn_bits_wdata [27] ), .QN(\EXU/_1304_ ) );
DFF_X1 \EXU/_2488_ ( .D(\EXU/_1556_ ), .CK(clock ), .Q(\_EXU_io_LSUIn_bits_wdata [28] ), .QN(\EXU/_1303_ ) );
DFF_X1 \EXU/_2489_ ( .D(\EXU/_1557_ ), .CK(clock ), .Q(\_EXU_io_LSUIn_bits_wdata [29] ), .QN(\EXU/_1302_ ) );
DFF_X1 \EXU/_2490_ ( .D(\EXU/_1558_ ), .CK(clock ), .Q(\_EXU_io_LSUIn_bits_wdata [30] ), .QN(\EXU/_1301_ ) );
DFF_X1 \EXU/_2491_ ( .D(\EXU/_1559_ ), .CK(clock ), .Q(\_EXU_io_LSUIn_bits_wdata [31] ), .QN(\EXU/_1300_ ) );
DFF_X1 \EXU/_2492_ ( .D(\EXU/_1560_ ), .CK(clock ), .Q(\EXU/in_imm [0] ), .QN(\EXU/_1299_ ) );
DFF_X1 \EXU/_2493_ ( .D(\EXU/_1561_ ), .CK(clock ), .Q(\EXU/in_imm [1] ), .QN(\EXU/_1298_ ) );
DFF_X1 \EXU/_2494_ ( .D(\EXU/_1562_ ), .CK(clock ), .Q(\EXU/in_imm [2] ), .QN(\EXU/_1297_ ) );
DFF_X1 \EXU/_2495_ ( .D(\EXU/_1563_ ), .CK(clock ), .Q(\EXU/in_imm [3] ), .QN(\EXU/_1296_ ) );
DFF_X1 \EXU/_2496_ ( .D(\EXU/_1564_ ), .CK(clock ), .Q(\EXU/in_imm [4] ), .QN(\EXU/_1295_ ) );
DFF_X1 \EXU/_2497_ ( .D(\EXU/_1565_ ), .CK(clock ), .Q(\EXU/in_imm [5] ), .QN(\EXU/_1294_ ) );
DFF_X1 \EXU/_2498_ ( .D(\EXU/_1566_ ), .CK(clock ), .Q(\EXU/in_imm [6] ), .QN(\EXU/_1293_ ) );
DFF_X1 \EXU/_2499_ ( .D(\EXU/_1567_ ), .CK(clock ), .Q(\EXU/in_imm [7] ), .QN(\EXU/_1292_ ) );
DFF_X1 \EXU/_2500_ ( .D(\EXU/_1568_ ), .CK(clock ), .Q(\EXU/in_imm [8] ), .QN(\EXU/_1291_ ) );
DFF_X1 \EXU/_2501_ ( .D(\EXU/_1569_ ), .CK(clock ), .Q(\EXU/in_imm [9] ), .QN(\EXU/_1290_ ) );
DFF_X1 \EXU/_2502_ ( .D(\EXU/_1570_ ), .CK(clock ), .Q(\EXU/in_imm [10] ), .QN(\EXU/_1289_ ) );
DFF_X1 \EXU/_2503_ ( .D(\EXU/_1571_ ), .CK(clock ), .Q(\EXU/in_imm [11] ), .QN(\EXU/_1288_ ) );
DFF_X1 \EXU/_2504_ ( .D(\EXU/_1572_ ), .CK(clock ), .Q(\EXU/in_imm [12] ), .QN(\EXU/_1287_ ) );
DFF_X1 \EXU/_2505_ ( .D(\EXU/_1573_ ), .CK(clock ), .Q(\EXU/in_imm [13] ), .QN(\EXU/_1286_ ) );
DFF_X1 \EXU/_2506_ ( .D(\EXU/_1574_ ), .CK(clock ), .Q(\EXU/in_imm [14] ), .QN(\EXU/_1285_ ) );
DFF_X1 \EXU/_2507_ ( .D(\EXU/_1575_ ), .CK(clock ), .Q(\EXU/in_imm [15] ), .QN(\EXU/_1284_ ) );
DFF_X1 \EXU/_2508_ ( .D(\EXU/_1576_ ), .CK(clock ), .Q(\EXU/in_imm [16] ), .QN(\EXU/_1283_ ) );
DFF_X1 \EXU/_2509_ ( .D(\EXU/_1577_ ), .CK(clock ), .Q(\EXU/in_imm [17] ), .QN(\EXU/_1282_ ) );
DFF_X1 \EXU/_2510_ ( .D(\EXU/_1578_ ), .CK(clock ), .Q(\EXU/in_imm [18] ), .QN(\EXU/_1281_ ) );
DFF_X1 \EXU/_2511_ ( .D(\EXU/_1579_ ), .CK(clock ), .Q(\EXU/in_imm [19] ), .QN(\EXU/_1280_ ) );
DFF_X1 \EXU/_2512_ ( .D(\EXU/_1580_ ), .CK(clock ), .Q(\EXU/in_imm [20] ), .QN(\EXU/_1279_ ) );
DFF_X1 \EXU/_2513_ ( .D(\EXU/_1581_ ), .CK(clock ), .Q(\EXU/in_imm [21] ), .QN(\EXU/_1278_ ) );
DFF_X1 \EXU/_2514_ ( .D(\EXU/_1582_ ), .CK(clock ), .Q(\EXU/in_imm [22] ), .QN(\EXU/_1277_ ) );
DFF_X1 \EXU/_2515_ ( .D(\EXU/_1583_ ), .CK(clock ), .Q(\EXU/in_imm [23] ), .QN(\EXU/_1276_ ) );
DFF_X1 \EXU/_2516_ ( .D(\EXU/_1584_ ), .CK(clock ), .Q(\EXU/in_imm [24] ), .QN(\EXU/_1275_ ) );
DFF_X1 \EXU/_2517_ ( .D(\EXU/_1585_ ), .CK(clock ), .Q(\EXU/in_imm [25] ), .QN(\EXU/_1274_ ) );
DFF_X1 \EXU/_2518_ ( .D(\EXU/_1586_ ), .CK(clock ), .Q(\EXU/in_imm [26] ), .QN(\EXU/_1273_ ) );
DFF_X1 \EXU/_2519_ ( .D(\EXU/_1587_ ), .CK(clock ), .Q(\EXU/in_imm [27] ), .QN(\EXU/_1272_ ) );
DFF_X1 \EXU/_2520_ ( .D(\EXU/_1588_ ), .CK(clock ), .Q(\EXU/in_imm [28] ), .QN(\EXU/_1271_ ) );
DFF_X1 \EXU/_2521_ ( .D(\EXU/_1589_ ), .CK(clock ), .Q(\EXU/in_imm [29] ), .QN(\EXU/_1270_ ) );
DFF_X1 \EXU/_2522_ ( .D(\EXU/_1590_ ), .CK(clock ), .Q(\EXU/in_imm [30] ), .QN(\EXU/_1269_ ) );
DFF_X1 \EXU/_2523_ ( .D(\EXU/_1591_ ), .CK(clock ), .Q(\EXU/in_imm [31] ), .QN(\EXU/_1268_ ) );
DFF_X1 \EXU/_2524_ ( .D(\EXU/_1592_ ), .CK(clock ), .Q(\EXU/in_uimm [0] ), .QN(\EXU/_1267_ ) );
DFF_X1 \EXU/_2525_ ( .D(\EXU/_1593_ ), .CK(clock ), .Q(\EXU/in_uimm [1] ), .QN(\EXU/_1266_ ) );
DFF_X1 \EXU/_2526_ ( .D(\EXU/_1594_ ), .CK(clock ), .Q(\EXU/in_uimm [2] ), .QN(\EXU/_1265_ ) );
DFF_X1 \EXU/_2527_ ( .D(\EXU/_1595_ ), .CK(clock ), .Q(\EXU/in_uimm [3] ), .QN(\EXU/_1264_ ) );
DFF_X1 \EXU/_2528_ ( .D(\EXU/_1596_ ), .CK(clock ), .Q(\EXU/in_uimm [4] ), .QN(\EXU/_1263_ ) );
DFF_X1 \EXU/_2529_ ( .D(\EXU/_1597_ ), .CK(clock ), .Q(\EXU/in_uimm [5] ), .QN(\EXU/_1262_ ) );
DFF_X1 \EXU/_2530_ ( .D(\EXU/_1598_ ), .CK(clock ), .Q(\EXU/in_uimm [6] ), .QN(\EXU/_1261_ ) );
DFF_X1 \EXU/_2531_ ( .D(\EXU/_1599_ ), .CK(clock ), .Q(\EXU/in_uimm [7] ), .QN(\EXU/_1260_ ) );
DFF_X1 \EXU/_2532_ ( .D(\EXU/_1600_ ), .CK(clock ), .Q(\EXU/in_uimm [8] ), .QN(\EXU/_1259_ ) );
DFF_X1 \EXU/_2533_ ( .D(\EXU/_1601_ ), .CK(clock ), .Q(\EXU/in_uimm [9] ), .QN(\EXU/_1258_ ) );
DFF_X1 \EXU/_2534_ ( .D(\EXU/_1602_ ), .CK(clock ), .Q(\EXU/in_uimm [10] ), .QN(\EXU/_1257_ ) );
DFF_X1 \EXU/_2535_ ( .D(\EXU/_1603_ ), .CK(clock ), .Q(\EXU/in_uimm [11] ), .QN(\EXU/_1256_ ) );
DFF_X1 \EXU/_2536_ ( .D(\EXU/_1604_ ), .CK(clock ), .Q(\EXU/in_uimm [12] ), .QN(\EXU/_1255_ ) );
DFF_X1 \EXU/_2537_ ( .D(\EXU/_1605_ ), .CK(clock ), .Q(\EXU/in_uimm [13] ), .QN(\EXU/_1254_ ) );
DFF_X1 \EXU/_2538_ ( .D(\EXU/_1606_ ), .CK(clock ), .Q(\EXU/in_uimm [14] ), .QN(\EXU/_1253_ ) );
DFF_X1 \EXU/_2539_ ( .D(\EXU/_1607_ ), .CK(clock ), .Q(\EXU/in_uimm [15] ), .QN(\EXU/_1252_ ) );
DFF_X1 \EXU/_2540_ ( .D(\EXU/_1608_ ), .CK(clock ), .Q(\EXU/in_uimm [16] ), .QN(\EXU/_1251_ ) );
DFF_X1 \EXU/_2541_ ( .D(\EXU/_1609_ ), .CK(clock ), .Q(\EXU/in_uimm [17] ), .QN(\EXU/_1250_ ) );
DFF_X1 \EXU/_2542_ ( .D(\EXU/_1610_ ), .CK(clock ), .Q(\EXU/in_uimm [18] ), .QN(\EXU/_1249_ ) );
DFF_X1 \EXU/_2543_ ( .D(\EXU/_1611_ ), .CK(clock ), .Q(\EXU/in_uimm [19] ), .QN(\EXU/_1248_ ) );
DFF_X1 \EXU/_2544_ ( .D(\EXU/_1612_ ), .CK(clock ), .Q(\EXU/in_uimm [20] ), .QN(\EXU/_1247_ ) );
DFF_X1 \EXU/_2545_ ( .D(\EXU/_1613_ ), .CK(clock ), .Q(\EXU/in_uimm [21] ), .QN(\EXU/_1246_ ) );
DFF_X1 \EXU/_2546_ ( .D(\EXU/_1614_ ), .CK(clock ), .Q(\EXU/in_uimm [22] ), .QN(\EXU/_1245_ ) );
DFF_X1 \EXU/_2547_ ( .D(\EXU/_1615_ ), .CK(clock ), .Q(\EXU/in_uimm [23] ), .QN(\EXU/_1244_ ) );
DFF_X1 \EXU/_2548_ ( .D(\EXU/_1616_ ), .CK(clock ), .Q(\EXU/in_uimm [24] ), .QN(\EXU/_1243_ ) );
DFF_X1 \EXU/_2549_ ( .D(\EXU/_1617_ ), .CK(clock ), .Q(\EXU/in_uimm [25] ), .QN(\EXU/_1242_ ) );
DFF_X1 \EXU/_2550_ ( .D(\EXU/_1618_ ), .CK(clock ), .Q(\EXU/in_uimm [26] ), .QN(\EXU/_1241_ ) );
DFF_X1 \EXU/_2551_ ( .D(\EXU/_1619_ ), .CK(clock ), .Q(\EXU/in_uimm [27] ), .QN(\EXU/_1240_ ) );
DFF_X1 \EXU/_2552_ ( .D(\EXU/_1620_ ), .CK(clock ), .Q(\EXU/in_uimm [28] ), .QN(\EXU/_1239_ ) );
DFF_X1 \EXU/_2553_ ( .D(\EXU/_1621_ ), .CK(clock ), .Q(\EXU/in_uimm [29] ), .QN(\EXU/_1238_ ) );
DFF_X1 \EXU/_2554_ ( .D(\EXU/_1622_ ), .CK(clock ), .Q(\EXU/in_uimm [30] ), .QN(\EXU/_1237_ ) );
DFF_X1 \EXU/_2555_ ( .D(\EXU/_1623_ ), .CK(clock ), .Q(\EXU/in_uimm [31] ), .QN(\EXU/_1236_ ) );
DFF_X1 \EXU/_2556_ ( .D(\EXU/_1624_ ), .CK(clock ), .Q(\EXU/in_control_aluASrc ), .QN(\EXU/_1235_ ) );
DFF_X1 \EXU/_2557_ ( .D(\EXU/_1625_ ), .CK(clock ), .Q(\EXU/in_control_aluBSrc [0] ), .QN(\EXU/_1234_ ) );
DFF_X1 \EXU/_2558_ ( .D(\EXU/_1626_ ), .CK(clock ), .Q(\EXU/in_control_aluBSrc [1] ), .QN(\EXU/_1233_ ) );
DFF_X1 \EXU/_2559_ ( .D(\EXU/_1627_ ), .CK(clock ), .Q(\EXU/in_control_aluCtr [0] ), .QN(\EXU/_1232_ ) );
DFF_X1 \EXU/_2560_ ( .D(\EXU/_1628_ ), .CK(clock ), .Q(\EXU/in_control_aluCtr [1] ), .QN(\EXU/_1231_ ) );
DFF_X1 \EXU/_2561_ ( .D(\EXU/_1629_ ), .CK(clock ), .Q(\EXU/in_control_aluCtr [2] ), .QN(\EXU/_1230_ ) );
DFF_X1 \EXU/_2562_ ( .D(\EXU/_1630_ ), .CK(clock ), .Q(\EXU/in_control_aluCtr [3] ), .QN(\EXU/_1229_ ) );
DFF_X1 \EXU/_2563_ ( .D(\EXU/_1631_ ), .CK(clock ), .Q(\EXU/in_control_csrSrc ), .QN(\EXU/_1228_ ) );
DFF_X1 \EXU/_2564_ ( .D(\EXU/_1632_ ), .CK(clock ), .Q(\EXU/in_control_csrCtr [0] ), .QN(\EXU/_1227_ ) );
DFF_X1 \EXU/_2565_ ( .D(\EXU/_1633_ ), .CK(clock ), .Q(\EXU/in_control_csrCtr [1] ), .QN(\EXU/_1226_ ) );
DFF_X1 \EXU/_2566_ ( .D(\EXU/_1634_ ), .CK(clock ), .Q(\EXU/in_control_csrCtr [2] ), .QN(\EXU/_1225_ ) );
DFF_X1 \EXU/_2567_ ( .D(\EXU/_1635_ ), .CK(clock ), .Q(\EXU/in_control_brType [0] ), .QN(\EXU/_1224_ ) );
DFF_X1 \EXU/_2568_ ( .D(\EXU/_1636_ ), .CK(clock ), .Q(\EXU/in_control_brType [1] ), .QN(\EXU/_1223_ ) );
DFF_X1 \EXU/_2569_ ( .D(\EXU/_1637_ ), .CK(clock ), .Q(\EXU/in_control_brType [2] ), .QN(\EXU/_1222_ ) );
DFF_X1 \EXU/_2570_ ( .D(\EXU/_1638_ ), .CK(clock ), .Q(_EXU_io_LSUIn_bits_ren ), .QN(\EXU/_1221_ ) );
DFF_X1 \EXU/_2571_ ( .D(\EXU/_1639_ ), .CK(clock ), .Q(_EXU_io_LSUIn_bits_wen ), .QN(\EXU/_1220_ ) );
DFF_X1 \EXU/_2572_ ( .D(\EXU/_1640_ ), .CK(clock ), .Q(\_EXU_io_LSUIn_bits_memOp [0] ), .QN(\EXU/_1219_ ) );
DFF_X1 \EXU/_2573_ ( .D(\EXU/_1641_ ), .CK(clock ), .Q(\_EXU_io_LSUIn_bits_memOp [1] ), .QN(\EXU/_1218_ ) );
DFF_X1 \EXU/_2574_ ( .D(\EXU/_1642_ ), .CK(clock ), .Q(\_EXU_io_LSUIn_bits_memOp [2] ), .QN(\EXU/_1217_ ) );
BUF_X1 \EXU/_2575_ ( .A(\_EXU_io_LSUIn_bits_raddr [0] ), .Z(\_EXU_io_LSUIn_bits_waddr [0] ) );
BUF_X1 \EXU/_2576_ ( .A(\_EXU_io_LSUIn_bits_raddr [1] ), .Z(\_EXU_io_LSUIn_bits_waddr [1] ) );
BUF_X1 \EXU/_2577_ ( .A(\_EXU_io_LSUIn_bits_raddr [2] ), .Z(\_EXU_io_LSUIn_bits_waddr [2] ) );
BUF_X1 \EXU/_2578_ ( .A(\_EXU_io_LSUIn_bits_raddr [3] ), .Z(\_EXU_io_LSUIn_bits_waddr [3] ) );
BUF_X1 \EXU/_2579_ ( .A(\_EXU_io_LSUIn_bits_raddr [4] ), .Z(\_EXU_io_LSUIn_bits_waddr [4] ) );
BUF_X1 \EXU/_2580_ ( .A(\_EXU_io_LSUIn_bits_raddr [5] ), .Z(\_EXU_io_LSUIn_bits_waddr [5] ) );
BUF_X1 \EXU/_2581_ ( .A(\_EXU_io_LSUIn_bits_raddr [6] ), .Z(\_EXU_io_LSUIn_bits_waddr [6] ) );
BUF_X1 \EXU/_2582_ ( .A(\_EXU_io_LSUIn_bits_raddr [7] ), .Z(\_EXU_io_LSUIn_bits_waddr [7] ) );
BUF_X1 \EXU/_2583_ ( .A(\_EXU_io_LSUIn_bits_raddr [8] ), .Z(\_EXU_io_LSUIn_bits_waddr [8] ) );
BUF_X1 \EXU/_2584_ ( .A(\_EXU_io_LSUIn_bits_raddr [9] ), .Z(\_EXU_io_LSUIn_bits_waddr [9] ) );
BUF_X1 \EXU/_2585_ ( .A(\_EXU_io_LSUIn_bits_raddr [10] ), .Z(\_EXU_io_LSUIn_bits_waddr [10] ) );
BUF_X1 \EXU/_2586_ ( .A(\_EXU_io_LSUIn_bits_raddr [11] ), .Z(\_EXU_io_LSUIn_bits_waddr [11] ) );
BUF_X1 \EXU/_2587_ ( .A(\_EXU_io_LSUIn_bits_raddr [12] ), .Z(\_EXU_io_LSUIn_bits_waddr [12] ) );
BUF_X1 \EXU/_2588_ ( .A(\_EXU_io_LSUIn_bits_raddr [13] ), .Z(\_EXU_io_LSUIn_bits_waddr [13] ) );
BUF_X1 \EXU/_2589_ ( .A(\_EXU_io_LSUIn_bits_raddr [14] ), .Z(\_EXU_io_LSUIn_bits_waddr [14] ) );
BUF_X1 \EXU/_2590_ ( .A(\_EXU_io_LSUIn_bits_raddr [15] ), .Z(\_EXU_io_LSUIn_bits_waddr [15] ) );
BUF_X1 \EXU/_2591_ ( .A(\_EXU_io_LSUIn_bits_raddr [16] ), .Z(\_EXU_io_LSUIn_bits_waddr [16] ) );
BUF_X1 \EXU/_2592_ ( .A(\_EXU_io_LSUIn_bits_raddr [17] ), .Z(\_EXU_io_LSUIn_bits_waddr [17] ) );
BUF_X1 \EXU/_2593_ ( .A(\_EXU_io_LSUIn_bits_raddr [18] ), .Z(\_EXU_io_LSUIn_bits_waddr [18] ) );
BUF_X1 \EXU/_2594_ ( .A(\_EXU_io_LSUIn_bits_raddr [19] ), .Z(\_EXU_io_LSUIn_bits_waddr [19] ) );
BUF_X1 \EXU/_2595_ ( .A(\_EXU_io_LSUIn_bits_raddr [20] ), .Z(\_EXU_io_LSUIn_bits_waddr [20] ) );
BUF_X1 \EXU/_2596_ ( .A(\_EXU_io_LSUIn_bits_raddr [21] ), .Z(\_EXU_io_LSUIn_bits_waddr [21] ) );
BUF_X1 \EXU/_2597_ ( .A(\_EXU_io_LSUIn_bits_raddr [22] ), .Z(\_EXU_io_LSUIn_bits_waddr [22] ) );
BUF_X1 \EXU/_2598_ ( .A(\_EXU_io_LSUIn_bits_raddr [23] ), .Z(\_EXU_io_LSUIn_bits_waddr [23] ) );
BUF_X1 \EXU/_2599_ ( .A(\_EXU_io_LSUIn_bits_raddr [24] ), .Z(\_EXU_io_LSUIn_bits_waddr [24] ) );
BUF_X1 \EXU/_2600_ ( .A(\_EXU_io_LSUIn_bits_raddr [25] ), .Z(\_EXU_io_LSUIn_bits_waddr [25] ) );
BUF_X1 \EXU/_2601_ ( .A(\_EXU_io_LSUIn_bits_raddr [26] ), .Z(\_EXU_io_LSUIn_bits_waddr [26] ) );
BUF_X1 \EXU/_2602_ ( .A(\_EXU_io_LSUIn_bits_raddr [27] ), .Z(\_EXU_io_LSUIn_bits_waddr [27] ) );
BUF_X1 \EXU/_2603_ ( .A(\_EXU_io_LSUIn_bits_raddr [28] ), .Z(\_EXU_io_LSUIn_bits_waddr [28] ) );
BUF_X1 \EXU/_2604_ ( .A(\_EXU_io_LSUIn_bits_raddr [29] ), .Z(\_EXU_io_LSUIn_bits_waddr [29] ) );
BUF_X1 \EXU/_2605_ ( .A(\_EXU_io_LSUIn_bits_raddr [30] ), .Z(\_EXU_io_LSUIn_bits_waddr [30] ) );
BUF_X1 \EXU/_2606_ ( .A(\_EXU_io_LSUIn_bits_raddr [31] ), .Z(\_EXU_io_LSUIn_bits_waddr [31] ) );
BUF_X1 \EXU/_2607_ ( .A(\_EXU_io_LSUIn_bits_raddr [0] ), .Z(\_EXU_io_out_bits_aluOut [0] ) );
BUF_X1 \EXU/_2608_ ( .A(\_EXU_io_LSUIn_bits_raddr [1] ), .Z(\_EXU_io_out_bits_aluOut [1] ) );
BUF_X1 \EXU/_2609_ ( .A(\_EXU_io_LSUIn_bits_raddr [2] ), .Z(\_EXU_io_out_bits_aluOut [2] ) );
BUF_X1 \EXU/_2610_ ( .A(\_EXU_io_LSUIn_bits_raddr [3] ), .Z(\_EXU_io_out_bits_aluOut [3] ) );
BUF_X1 \EXU/_2611_ ( .A(\_EXU_io_LSUIn_bits_raddr [4] ), .Z(\_EXU_io_out_bits_aluOut [4] ) );
BUF_X1 \EXU/_2612_ ( .A(\_EXU_io_LSUIn_bits_raddr [5] ), .Z(\_EXU_io_out_bits_aluOut [5] ) );
BUF_X1 \EXU/_2613_ ( .A(\_EXU_io_LSUIn_bits_raddr [6] ), .Z(\_EXU_io_out_bits_aluOut [6] ) );
BUF_X1 \EXU/_2614_ ( .A(\_EXU_io_LSUIn_bits_raddr [7] ), .Z(\_EXU_io_out_bits_aluOut [7] ) );
BUF_X1 \EXU/_2615_ ( .A(\_EXU_io_LSUIn_bits_raddr [8] ), .Z(\_EXU_io_out_bits_aluOut [8] ) );
BUF_X1 \EXU/_2616_ ( .A(\_EXU_io_LSUIn_bits_raddr [9] ), .Z(\_EXU_io_out_bits_aluOut [9] ) );
BUF_X1 \EXU/_2617_ ( .A(\_EXU_io_LSUIn_bits_raddr [10] ), .Z(\_EXU_io_out_bits_aluOut [10] ) );
BUF_X1 \EXU/_2618_ ( .A(\_EXU_io_LSUIn_bits_raddr [11] ), .Z(\_EXU_io_out_bits_aluOut [11] ) );
BUF_X1 \EXU/_2619_ ( .A(\_EXU_io_LSUIn_bits_raddr [12] ), .Z(\_EXU_io_out_bits_aluOut [12] ) );
BUF_X1 \EXU/_2620_ ( .A(\_EXU_io_LSUIn_bits_raddr [13] ), .Z(\_EXU_io_out_bits_aluOut [13] ) );
BUF_X1 \EXU/_2621_ ( .A(\_EXU_io_LSUIn_bits_raddr [14] ), .Z(\_EXU_io_out_bits_aluOut [14] ) );
BUF_X1 \EXU/_2622_ ( .A(\_EXU_io_LSUIn_bits_raddr [15] ), .Z(\_EXU_io_out_bits_aluOut [15] ) );
BUF_X1 \EXU/_2623_ ( .A(\_EXU_io_LSUIn_bits_raddr [16] ), .Z(\_EXU_io_out_bits_aluOut [16] ) );
BUF_X1 \EXU/_2624_ ( .A(\_EXU_io_LSUIn_bits_raddr [17] ), .Z(\_EXU_io_out_bits_aluOut [17] ) );
BUF_X1 \EXU/_2625_ ( .A(\_EXU_io_LSUIn_bits_raddr [18] ), .Z(\_EXU_io_out_bits_aluOut [18] ) );
BUF_X1 \EXU/_2626_ ( .A(\_EXU_io_LSUIn_bits_raddr [19] ), .Z(\_EXU_io_out_bits_aluOut [19] ) );
BUF_X1 \EXU/_2627_ ( .A(\_EXU_io_LSUIn_bits_raddr [20] ), .Z(\_EXU_io_out_bits_aluOut [20] ) );
BUF_X1 \EXU/_2628_ ( .A(\_EXU_io_LSUIn_bits_raddr [21] ), .Z(\_EXU_io_out_bits_aluOut [21] ) );
BUF_X1 \EXU/_2629_ ( .A(\_EXU_io_LSUIn_bits_raddr [22] ), .Z(\_EXU_io_out_bits_aluOut [22] ) );
BUF_X1 \EXU/_2630_ ( .A(\_EXU_io_LSUIn_bits_raddr [23] ), .Z(\_EXU_io_out_bits_aluOut [23] ) );
BUF_X1 \EXU/_2631_ ( .A(\_EXU_io_LSUIn_bits_raddr [24] ), .Z(\_EXU_io_out_bits_aluOut [24] ) );
BUF_X1 \EXU/_2632_ ( .A(\_EXU_io_LSUIn_bits_raddr [25] ), .Z(\_EXU_io_out_bits_aluOut [25] ) );
BUF_X1 \EXU/_2633_ ( .A(\_EXU_io_LSUIn_bits_raddr [26] ), .Z(\_EXU_io_out_bits_aluOut [26] ) );
BUF_X1 \EXU/_2634_ ( .A(\_EXU_io_LSUIn_bits_raddr [27] ), .Z(\_EXU_io_out_bits_aluOut [27] ) );
BUF_X1 \EXU/_2635_ ( .A(\_EXU_io_LSUIn_bits_raddr [28] ), .Z(\_EXU_io_out_bits_aluOut [28] ) );
BUF_X1 \EXU/_2636_ ( .A(\_EXU_io_LSUIn_bits_raddr [29] ), .Z(\_EXU_io_out_bits_aluOut [29] ) );
BUF_X1 \EXU/_2637_ ( .A(\_EXU_io_LSUIn_bits_raddr [30] ), .Z(\_EXU_io_out_bits_aluOut [30] ) );
BUF_X1 \EXU/_2638_ ( .A(\_EXU_io_LSUIn_bits_raddr [31] ), .Z(\_EXU_io_out_bits_aluOut [31] ) );
BUF_X1 \EXU/_2639_ ( .A(_IDU_io_out_bits_control_pcSrc ), .Z(_EXU_io_out_bits_control_pcSrc ) );
BUF_X1 \EXU/_2640_ ( .A(_IDU_io_out_bits_control_regWe ), .Z(_EXU_io_out_bits_control_regWe ) );
BUF_X1 \EXU/_2641_ ( .A(\_IDU_io_out_bits_control_wbSrc [0] ), .Z(\_EXU_io_out_bits_control_wbSrc [0] ) );
BUF_X1 \EXU/_2642_ ( .A(\_IDU_io_out_bits_control_wbSrc [1] ), .Z(\_EXU_io_out_bits_control_wbSrc [1] ) );
BUF_X1 \EXU/_2643_ ( .A(\_IDU_io_out_bits_wa [0] ), .Z(\_EXU_io_out_bits_wa [0] ) );
BUF_X1 \EXU/_2644_ ( .A(\_IDU_io_out_bits_wa [1] ), .Z(\_EXU_io_out_bits_wa [1] ) );
BUF_X1 \EXU/_2645_ ( .A(\_IDU_io_out_bits_wa [2] ), .Z(\_EXU_io_out_bits_wa [2] ) );
BUF_X1 \EXU/_2646_ ( .A(\_IDU_io_out_bits_wa [3] ), .Z(\_EXU_io_out_bits_wa [3] ) );
BUF_X1 \EXU/_2647_ ( .A(\_IDU_io_out_bits_wa [4] ), .Z(\_EXU_io_out_bits_wa [4] ) );
BUF_X1 \EXU/_2648_ ( .A(\EXU/state [0] ), .Z(\EXU/_1215_ ) );
BUF_X1 \EXU/_2649_ ( .A(\EXU/state [1] ), .Z(\EXU/_1216_ ) );
BUF_X1 \EXU/_2650_ ( .A(\EXU/_0842_ ), .Z(_EXU_io_out_valid ) );
BUF_X1 \EXU/_2651_ ( .A(\EXU/_0594_ ), .Z(_EXU_io_LSUOut_ready ) );
BUF_X1 \EXU/_2652_ ( .A(\EXU/_0561_ ), .Z(_EXU_io_LSUIn_valid ) );
BUF_X1 \EXU/_2653_ ( .A(\EXU/_0775_ ), .Z(_EXU_io_in_ready ) );
BUF_X1 \EXU/_2654_ ( .A(_IDU_io_out_valid ), .Z(\EXU/_0776_ ) );
BUF_X1 \EXU/_2655_ ( .A(\EXU/in_rd1 [0] ), .Z(\EXU/_0459_ ) );
BUF_X1 \EXU/_2656_ ( .A(\EXU/in_pc [0] ), .Z(\EXU/_0427_ ) );
BUF_X1 \EXU/_2657_ ( .A(\EXU/in_control_aluASrc ), .Z(\EXU/_0381_ ) );
BUF_X1 \EXU/_2658_ ( .A(\EXU/_0069_ ), .Z(\EXU/_0000_ ) );
BUF_X1 \EXU/_2659_ ( .A(\EXU/in_rd1 [1] ), .Z(\EXU/_0470_ ) );
BUF_X1 \EXU/_2660_ ( .A(\EXU/in_pc [1] ), .Z(\EXU/_0438_ ) );
BUF_X1 \EXU/_2661_ ( .A(\EXU/_0080_ ), .Z(\EXU/_0011_ ) );
BUF_X1 \EXU/_2662_ ( .A(\EXU/in_rd1 [2] ), .Z(\EXU/_0481_ ) );
BUF_X1 \EXU/_2663_ ( .A(\EXU/in_pc [2] ), .Z(\EXU/_0449_ ) );
BUF_X1 \EXU/_2664_ ( .A(\EXU/_0091_ ), .Z(\EXU/_0022_ ) );
BUF_X1 \EXU/_2665_ ( .A(\EXU/in_rd1 [3] ), .Z(\EXU/_0484_ ) );
BUF_X1 \EXU/_2666_ ( .A(\EXU/in_pc [3] ), .Z(\EXU/_0452_ ) );
BUF_X1 \EXU/_2667_ ( .A(\EXU/_0094_ ), .Z(\EXU/_0025_ ) );
BUF_X1 \EXU/_2668_ ( .A(\EXU/in_rd1 [4] ), .Z(\EXU/_0485_ ) );
BUF_X1 \EXU/_2669_ ( .A(\EXU/in_pc [4] ), .Z(\EXU/_0453_ ) );
BUF_X1 \EXU/_2670_ ( .A(\EXU/_0095_ ), .Z(\EXU/_0026_ ) );
BUF_X1 \EXU/_2671_ ( .A(\EXU/in_rd1 [5] ), .Z(\EXU/_0486_ ) );
BUF_X1 \EXU/_2672_ ( .A(\EXU/in_pc [5] ), .Z(\EXU/_0454_ ) );
BUF_X1 \EXU/_2673_ ( .A(\EXU/_0096_ ), .Z(\EXU/_0027_ ) );
BUF_X1 \EXU/_2674_ ( .A(\EXU/in_rd1 [6] ), .Z(\EXU/_0487_ ) );
BUF_X1 \EXU/_2675_ ( .A(\EXU/in_pc [6] ), .Z(\EXU/_0455_ ) );
BUF_X1 \EXU/_2676_ ( .A(\EXU/_0097_ ), .Z(\EXU/_0028_ ) );
BUF_X1 \EXU/_2677_ ( .A(\EXU/in_rd1 [7] ), .Z(\EXU/_0488_ ) );
BUF_X1 \EXU/_2678_ ( .A(\EXU/in_pc [7] ), .Z(\EXU/_0456_ ) );
BUF_X1 \EXU/_2679_ ( .A(\EXU/_0098_ ), .Z(\EXU/_0029_ ) );
BUF_X1 \EXU/_2680_ ( .A(\EXU/in_rd1 [8] ), .Z(\EXU/_0489_ ) );
BUF_X1 \EXU/_2681_ ( .A(\EXU/in_pc [8] ), .Z(\EXU/_0457_ ) );
BUF_X1 \EXU/_2682_ ( .A(\EXU/_0099_ ), .Z(\EXU/_0030_ ) );
BUF_X1 \EXU/_2683_ ( .A(\EXU/in_rd1 [9] ), .Z(\EXU/_0490_ ) );
BUF_X1 \EXU/_2684_ ( .A(\EXU/in_pc [9] ), .Z(\EXU/_0458_ ) );
BUF_X1 \EXU/_2685_ ( .A(\EXU/_0100_ ), .Z(\EXU/_0031_ ) );
BUF_X1 \EXU/_2686_ ( .A(\EXU/in_rd1 [10] ), .Z(\EXU/_0460_ ) );
BUF_X1 \EXU/_2687_ ( .A(\EXU/in_pc [10] ), .Z(\EXU/_0428_ ) );
BUF_X1 \EXU/_2688_ ( .A(\EXU/_0070_ ), .Z(\EXU/_0001_ ) );
BUF_X1 \EXU/_2689_ ( .A(\EXU/in_rd1 [11] ), .Z(\EXU/_0461_ ) );
BUF_X1 \EXU/_2690_ ( .A(\EXU/in_pc [11] ), .Z(\EXU/_0429_ ) );
BUF_X1 \EXU/_2691_ ( .A(\EXU/_0071_ ), .Z(\EXU/_0002_ ) );
BUF_X1 \EXU/_2692_ ( .A(\EXU/in_rd1 [12] ), .Z(\EXU/_0462_ ) );
BUF_X1 \EXU/_2693_ ( .A(\EXU/in_pc [12] ), .Z(\EXU/_0430_ ) );
BUF_X1 \EXU/_2694_ ( .A(\EXU/_0072_ ), .Z(\EXU/_0003_ ) );
BUF_X1 \EXU/_2695_ ( .A(\EXU/in_rd1 [13] ), .Z(\EXU/_0463_ ) );
BUF_X1 \EXU/_2696_ ( .A(\EXU/in_pc [13] ), .Z(\EXU/_0431_ ) );
BUF_X1 \EXU/_2697_ ( .A(\EXU/_0073_ ), .Z(\EXU/_0004_ ) );
BUF_X1 \EXU/_2698_ ( .A(\EXU/in_rd1 [14] ), .Z(\EXU/_0464_ ) );
BUF_X1 \EXU/_2699_ ( .A(\EXU/in_pc [14] ), .Z(\EXU/_0432_ ) );
BUF_X1 \EXU/_2700_ ( .A(\EXU/_0074_ ), .Z(\EXU/_0005_ ) );
BUF_X1 \EXU/_2701_ ( .A(\EXU/in_rd1 [15] ), .Z(\EXU/_0465_ ) );
BUF_X1 \EXU/_2702_ ( .A(\EXU/in_pc [15] ), .Z(\EXU/_0433_ ) );
BUF_X1 \EXU/_2703_ ( .A(\EXU/_0075_ ), .Z(\EXU/_0006_ ) );
BUF_X1 \EXU/_2704_ ( .A(\EXU/in_rd1 [16] ), .Z(\EXU/_0466_ ) );
BUF_X1 \EXU/_2705_ ( .A(\EXU/in_pc [16] ), .Z(\EXU/_0434_ ) );
BUF_X1 \EXU/_2706_ ( .A(\EXU/_0076_ ), .Z(\EXU/_0007_ ) );
BUF_X1 \EXU/_2707_ ( .A(\EXU/in_rd1 [17] ), .Z(\EXU/_0467_ ) );
BUF_X1 \EXU/_2708_ ( .A(\EXU/in_pc [17] ), .Z(\EXU/_0435_ ) );
BUF_X1 \EXU/_2709_ ( .A(\EXU/_0077_ ), .Z(\EXU/_0008_ ) );
BUF_X1 \EXU/_2710_ ( .A(\EXU/in_rd1 [18] ), .Z(\EXU/_0468_ ) );
BUF_X1 \EXU/_2711_ ( .A(\EXU/in_pc [18] ), .Z(\EXU/_0436_ ) );
BUF_X1 \EXU/_2712_ ( .A(\EXU/_0078_ ), .Z(\EXU/_0009_ ) );
BUF_X1 \EXU/_2713_ ( .A(\EXU/in_rd1 [19] ), .Z(\EXU/_0469_ ) );
BUF_X1 \EXU/_2714_ ( .A(\EXU/in_pc [19] ), .Z(\EXU/_0437_ ) );
BUF_X1 \EXU/_2715_ ( .A(\EXU/_0079_ ), .Z(\EXU/_0010_ ) );
BUF_X1 \EXU/_2716_ ( .A(\EXU/in_rd1 [20] ), .Z(\EXU/_0471_ ) );
BUF_X1 \EXU/_2717_ ( .A(\EXU/in_pc [20] ), .Z(\EXU/_0439_ ) );
BUF_X1 \EXU/_2718_ ( .A(\EXU/_0081_ ), .Z(\EXU/_0012_ ) );
BUF_X1 \EXU/_2719_ ( .A(\EXU/in_rd1 [21] ), .Z(\EXU/_0472_ ) );
BUF_X1 \EXU/_2720_ ( .A(\EXU/in_pc [21] ), .Z(\EXU/_0440_ ) );
BUF_X1 \EXU/_2721_ ( .A(\EXU/_0082_ ), .Z(\EXU/_0013_ ) );
BUF_X1 \EXU/_2722_ ( .A(\EXU/in_rd1 [22] ), .Z(\EXU/_0473_ ) );
BUF_X1 \EXU/_2723_ ( .A(\EXU/in_pc [22] ), .Z(\EXU/_0441_ ) );
BUF_X1 \EXU/_2724_ ( .A(\EXU/_0083_ ), .Z(\EXU/_0014_ ) );
BUF_X1 \EXU/_2725_ ( .A(\EXU/in_rd1 [23] ), .Z(\EXU/_0474_ ) );
BUF_X1 \EXU/_2726_ ( .A(\EXU/in_pc [23] ), .Z(\EXU/_0442_ ) );
BUF_X1 \EXU/_2727_ ( .A(\EXU/_0084_ ), .Z(\EXU/_0015_ ) );
BUF_X1 \EXU/_2728_ ( .A(\EXU/in_rd1 [24] ), .Z(\EXU/_0475_ ) );
BUF_X1 \EXU/_2729_ ( .A(\EXU/in_pc [24] ), .Z(\EXU/_0443_ ) );
BUF_X1 \EXU/_2730_ ( .A(\EXU/_0085_ ), .Z(\EXU/_0016_ ) );
BUF_X1 \EXU/_2731_ ( .A(\EXU/in_rd1 [25] ), .Z(\EXU/_0476_ ) );
BUF_X1 \EXU/_2732_ ( .A(\EXU/in_pc [25] ), .Z(\EXU/_0444_ ) );
BUF_X1 \EXU/_2733_ ( .A(\EXU/_0086_ ), .Z(\EXU/_0017_ ) );
BUF_X1 \EXU/_2734_ ( .A(\EXU/in_rd1 [26] ), .Z(\EXU/_0477_ ) );
BUF_X1 \EXU/_2735_ ( .A(\EXU/in_pc [26] ), .Z(\EXU/_0445_ ) );
BUF_X1 \EXU/_2736_ ( .A(\EXU/_0087_ ), .Z(\EXU/_0018_ ) );
BUF_X1 \EXU/_2737_ ( .A(\EXU/in_rd1 [27] ), .Z(\EXU/_0478_ ) );
BUF_X1 \EXU/_2738_ ( .A(\EXU/in_pc [27] ), .Z(\EXU/_0446_ ) );
BUF_X1 \EXU/_2739_ ( .A(\EXU/_0088_ ), .Z(\EXU/_0019_ ) );
BUF_X1 \EXU/_2740_ ( .A(\EXU/in_rd1 [28] ), .Z(\EXU/_0479_ ) );
BUF_X1 \EXU/_2741_ ( .A(\EXU/in_pc [28] ), .Z(\EXU/_0447_ ) );
BUF_X1 \EXU/_2742_ ( .A(\EXU/_0089_ ), .Z(\EXU/_0020_ ) );
BUF_X1 \EXU/_2743_ ( .A(\EXU/in_rd1 [29] ), .Z(\EXU/_0480_ ) );
BUF_X1 \EXU/_2744_ ( .A(\EXU/in_pc [29] ), .Z(\EXU/_0448_ ) );
BUF_X1 \EXU/_2745_ ( .A(\EXU/_0090_ ), .Z(\EXU/_0021_ ) );
BUF_X1 \EXU/_2746_ ( .A(\EXU/in_rd1 [30] ), .Z(\EXU/_0482_ ) );
BUF_X1 \EXU/_2747_ ( .A(\EXU/in_pc [30] ), .Z(\EXU/_0450_ ) );
BUF_X1 \EXU/_2748_ ( .A(\EXU/_0092_ ), .Z(\EXU/_0023_ ) );
BUF_X1 \EXU/_2749_ ( .A(\EXU/in_rd1 [31] ), .Z(\EXU/_0483_ ) );
BUF_X1 \EXU/_2750_ ( .A(\EXU/in_pc [31] ), .Z(\EXU/_0451_ ) );
BUF_X1 \EXU/_2751_ ( .A(\EXU/_0093_ ), .Z(\EXU/_0024_ ) );
BUF_X1 \EXU/_2752_ ( .A(\EXU/in_control_csrCtr [0] ), .Z(\EXU/_0391_ ) );
BUF_X1 \EXU/_2753_ ( .A(\EXU/_0101_ ), .Z(\EXU/_0032_ ) );
BUF_X1 \EXU/_2754_ ( .A(\EXU/in_control_csrCtr [1] ), .Z(\EXU/_0392_ ) );
BUF_X1 \EXU/_2755_ ( .A(\EXU/_0102_ ), .Z(\EXU/_0033_ ) );
BUF_X1 \EXU/_2756_ ( .A(\EXU/in_control_csrCtr [2] ), .Z(\EXU/_0393_ ) );
BUF_X1 \EXU/_2757_ ( .A(\EXU/_0103_ ), .Z(\EXU/_0034_ ) );
BUF_X1 \EXU/_2758_ ( .A(\EXU/in_uimm [0] ), .Z(\EXU/_0491_ ) );
BUF_X1 \EXU/_2759_ ( .A(\EXU/in_control_csrSrc ), .Z(\EXU/_0394_ ) );
BUF_X1 \EXU/_2760_ ( .A(\EXU/_0104_ ), .Z(\EXU/_0035_ ) );
BUF_X1 \EXU/_2761_ ( .A(\EXU/in_uimm [1] ), .Z(\EXU/_0502_ ) );
BUF_X1 \EXU/_2762_ ( .A(\EXU/_0115_ ), .Z(\EXU/_0046_ ) );
BUF_X1 \EXU/_2763_ ( .A(\EXU/in_uimm [2] ), .Z(\EXU/_0513_ ) );
BUF_X1 \EXU/_2764_ ( .A(\EXU/_0126_ ), .Z(\EXU/_0057_ ) );
BUF_X1 \EXU/_2765_ ( .A(\EXU/in_uimm [3] ), .Z(\EXU/_0516_ ) );
BUF_X1 \EXU/_2766_ ( .A(\EXU/_0129_ ), .Z(\EXU/_0060_ ) );
BUF_X1 \EXU/_2767_ ( .A(\EXU/in_uimm [4] ), .Z(\EXU/_0517_ ) );
BUF_X1 \EXU/_2768_ ( .A(\EXU/_0130_ ), .Z(\EXU/_0061_ ) );
BUF_X1 \EXU/_2769_ ( .A(\EXU/in_uimm [5] ), .Z(\EXU/_0518_ ) );
BUF_X1 \EXU/_2770_ ( .A(\EXU/_0131_ ), .Z(\EXU/_0062_ ) );
BUF_X1 \EXU/_2771_ ( .A(\EXU/in_uimm [6] ), .Z(\EXU/_0519_ ) );
BUF_X1 \EXU/_2772_ ( .A(\EXU/_0132_ ), .Z(\EXU/_0063_ ) );
BUF_X1 \EXU/_2773_ ( .A(\EXU/in_uimm [7] ), .Z(\EXU/_0520_ ) );
BUF_X1 \EXU/_2774_ ( .A(\EXU/_0133_ ), .Z(\EXU/_0064_ ) );
BUF_X1 \EXU/_2775_ ( .A(\EXU/in_uimm [8] ), .Z(\EXU/_0521_ ) );
BUF_X1 \EXU/_2776_ ( .A(\EXU/_0134_ ), .Z(\EXU/_0065_ ) );
BUF_X1 \EXU/_2777_ ( .A(\EXU/in_uimm [9] ), .Z(\EXU/_0522_ ) );
BUF_X1 \EXU/_2778_ ( .A(\EXU/_0135_ ), .Z(\EXU/_0066_ ) );
BUF_X1 \EXU/_2779_ ( .A(\EXU/in_uimm [10] ), .Z(\EXU/_0492_ ) );
BUF_X1 \EXU/_2780_ ( .A(\EXU/_0105_ ), .Z(\EXU/_0036_ ) );
BUF_X1 \EXU/_2781_ ( .A(\EXU/in_uimm [11] ), .Z(\EXU/_0493_ ) );
BUF_X1 \EXU/_2782_ ( .A(\EXU/_0106_ ), .Z(\EXU/_0037_ ) );
BUF_X1 \EXU/_2783_ ( .A(\EXU/in_uimm [12] ), .Z(\EXU/_0494_ ) );
BUF_X1 \EXU/_2784_ ( .A(\EXU/_0107_ ), .Z(\EXU/_0038_ ) );
BUF_X1 \EXU/_2785_ ( .A(\EXU/in_uimm [13] ), .Z(\EXU/_0495_ ) );
BUF_X1 \EXU/_2786_ ( .A(\EXU/_0108_ ), .Z(\EXU/_0039_ ) );
BUF_X1 \EXU/_2787_ ( .A(\EXU/in_uimm [14] ), .Z(\EXU/_0496_ ) );
BUF_X1 \EXU/_2788_ ( .A(\EXU/_0109_ ), .Z(\EXU/_0040_ ) );
BUF_X1 \EXU/_2789_ ( .A(\EXU/in_uimm [15] ), .Z(\EXU/_0497_ ) );
BUF_X1 \EXU/_2790_ ( .A(\EXU/_0110_ ), .Z(\EXU/_0041_ ) );
BUF_X1 \EXU/_2791_ ( .A(\EXU/in_uimm [16] ), .Z(\EXU/_0498_ ) );
BUF_X1 \EXU/_2792_ ( .A(\EXU/_0111_ ), .Z(\EXU/_0042_ ) );
BUF_X1 \EXU/_2793_ ( .A(\EXU/in_uimm [17] ), .Z(\EXU/_0499_ ) );
BUF_X1 \EXU/_2794_ ( .A(\EXU/_0112_ ), .Z(\EXU/_0043_ ) );
BUF_X1 \EXU/_2795_ ( .A(\EXU/in_uimm [18] ), .Z(\EXU/_0500_ ) );
BUF_X1 \EXU/_2796_ ( .A(\EXU/_0113_ ), .Z(\EXU/_0044_ ) );
BUF_X1 \EXU/_2797_ ( .A(\EXU/in_uimm [19] ), .Z(\EXU/_0501_ ) );
BUF_X1 \EXU/_2798_ ( .A(\EXU/_0114_ ), .Z(\EXU/_0045_ ) );
BUF_X1 \EXU/_2799_ ( .A(\EXU/in_uimm [20] ), .Z(\EXU/_0503_ ) );
BUF_X1 \EXU/_2800_ ( .A(\EXU/_0116_ ), .Z(\EXU/_0047_ ) );
BUF_X1 \EXU/_2801_ ( .A(\EXU/in_uimm [21] ), .Z(\EXU/_0504_ ) );
BUF_X1 \EXU/_2802_ ( .A(\EXU/_0117_ ), .Z(\EXU/_0048_ ) );
BUF_X1 \EXU/_2803_ ( .A(\EXU/in_uimm [22] ), .Z(\EXU/_0505_ ) );
BUF_X1 \EXU/_2804_ ( .A(\EXU/_0118_ ), .Z(\EXU/_0049_ ) );
BUF_X1 \EXU/_2805_ ( .A(\EXU/in_uimm [23] ), .Z(\EXU/_0506_ ) );
BUF_X1 \EXU/_2806_ ( .A(\EXU/_0119_ ), .Z(\EXU/_0050_ ) );
BUF_X1 \EXU/_2807_ ( .A(\EXU/in_uimm [24] ), .Z(\EXU/_0507_ ) );
BUF_X1 \EXU/_2808_ ( .A(\EXU/_0120_ ), .Z(\EXU/_0051_ ) );
BUF_X1 \EXU/_2809_ ( .A(\EXU/in_uimm [25] ), .Z(\EXU/_0508_ ) );
BUF_X1 \EXU/_2810_ ( .A(\EXU/_0121_ ), .Z(\EXU/_0052_ ) );
BUF_X1 \EXU/_2811_ ( .A(\EXU/in_uimm [26] ), .Z(\EXU/_0509_ ) );
BUF_X1 \EXU/_2812_ ( .A(\EXU/_0122_ ), .Z(\EXU/_0053_ ) );
BUF_X1 \EXU/_2813_ ( .A(\EXU/in_uimm [27] ), .Z(\EXU/_0510_ ) );
BUF_X1 \EXU/_2814_ ( .A(\EXU/_0123_ ), .Z(\EXU/_0054_ ) );
BUF_X1 \EXU/_2815_ ( .A(\EXU/in_uimm [28] ), .Z(\EXU/_0511_ ) );
BUF_X1 \EXU/_2816_ ( .A(\EXU/_0124_ ), .Z(\EXU/_0055_ ) );
BUF_X1 \EXU/_2817_ ( .A(\EXU/in_uimm [29] ), .Z(\EXU/_0512_ ) );
BUF_X1 \EXU/_2818_ ( .A(\EXU/_0125_ ), .Z(\EXU/_0056_ ) );
BUF_X1 \EXU/_2819_ ( .A(\EXU/in_uimm [30] ), .Z(\EXU/_0514_ ) );
BUF_X1 \EXU/_2820_ ( .A(\EXU/_0127_ ), .Z(\EXU/_0058_ ) );
BUF_X1 \EXU/_2821_ ( .A(\EXU/in_uimm [31] ), .Z(\EXU/_0515_ ) );
BUF_X1 \EXU/_2822_ ( .A(\EXU/_0128_ ), .Z(\EXU/_0059_ ) );
BUF_X1 \EXU/_2823_ ( .A(\EXU/in_control_aluBSrc [0] ), .Z(\EXU/_0382_ ) );
BUF_X1 \EXU/_2824_ ( .A(\EXU/in_control_aluBSrc [1] ), .Z(\EXU/_0383_ ) );
BUF_X1 \EXU/_2825_ ( .A(\EXU/in_imm [0] ), .Z(\EXU/_0395_ ) );
BUF_X1 \EXU/_2826_ ( .A(\_EXU_io_LSUIn_bits_wdata [0] ), .Z(\EXU/_0527_ ) );
BUF_X1 \EXU/_2827_ ( .A(\EXU/_0349_ ), .Z(\EXU/casez_tmp_0 [0] ) );
BUF_X1 \EXU/_2828_ ( .A(\EXU/in_imm [1] ), .Z(\EXU/_0406_ ) );
BUF_X1 \EXU/_2829_ ( .A(\_EXU_io_LSUIn_bits_wdata [1] ), .Z(\EXU/_0538_ ) );
BUF_X1 \EXU/_2830_ ( .A(\EXU/_0360_ ), .Z(\EXU/casez_tmp_0 [1] ) );
BUF_X1 \EXU/_2831_ ( .A(\EXU/in_imm [2] ), .Z(\EXU/_0417_ ) );
BUF_X1 \EXU/_2832_ ( .A(\_EXU_io_LSUIn_bits_wdata [2] ), .Z(\EXU/_0549_ ) );
BUF_X1 \EXU/_2833_ ( .A(\EXU/_0371_ ), .Z(\EXU/casez_tmp_0 [2] ) );
BUF_X1 \EXU/_2834_ ( .A(\EXU/in_imm [3] ), .Z(\EXU/_0420_ ) );
BUF_X1 \EXU/_2835_ ( .A(\_EXU_io_LSUIn_bits_wdata [3] ), .Z(\EXU/_0552_ ) );
BUF_X1 \EXU/_2836_ ( .A(\EXU/_0374_ ), .Z(\EXU/casez_tmp_0 [3] ) );
BUF_X1 \EXU/_2837_ ( .A(\EXU/in_imm [4] ), .Z(\EXU/_0421_ ) );
BUF_X1 \EXU/_2838_ ( .A(\_EXU_io_LSUIn_bits_wdata [4] ), .Z(\EXU/_0553_ ) );
BUF_X1 \EXU/_2839_ ( .A(\EXU/_0375_ ), .Z(\EXU/casez_tmp_0 [4] ) );
BUF_X1 \EXU/_2840_ ( .A(\EXU/in_imm [5] ), .Z(\EXU/_0422_ ) );
BUF_X1 \EXU/_2841_ ( .A(\_EXU_io_LSUIn_bits_wdata [5] ), .Z(\EXU/_0554_ ) );
BUF_X1 \EXU/_2842_ ( .A(\EXU/_0376_ ), .Z(\EXU/casez_tmp_0 [5] ) );
BUF_X1 \EXU/_2843_ ( .A(\EXU/in_imm [6] ), .Z(\EXU/_0423_ ) );
BUF_X1 \EXU/_2844_ ( .A(\_EXU_io_LSUIn_bits_wdata [6] ), .Z(\EXU/_0555_ ) );
BUF_X1 \EXU/_2845_ ( .A(\EXU/_0377_ ), .Z(\EXU/casez_tmp_0 [6] ) );
BUF_X1 \EXU/_2846_ ( .A(\EXU/in_imm [7] ), .Z(\EXU/_0424_ ) );
BUF_X1 \EXU/_2847_ ( .A(\_EXU_io_LSUIn_bits_wdata [7] ), .Z(\EXU/_0556_ ) );
BUF_X1 \EXU/_2848_ ( .A(\EXU/_0378_ ), .Z(\EXU/casez_tmp_0 [7] ) );
BUF_X1 \EXU/_2849_ ( .A(\EXU/in_imm [8] ), .Z(\EXU/_0425_ ) );
BUF_X1 \EXU/_2850_ ( .A(\_EXU_io_LSUIn_bits_wdata [8] ), .Z(\EXU/_0557_ ) );
BUF_X1 \EXU/_2851_ ( .A(\EXU/_0379_ ), .Z(\EXU/casez_tmp_0 [8] ) );
BUF_X1 \EXU/_2852_ ( .A(\EXU/in_imm [9] ), .Z(\EXU/_0426_ ) );
BUF_X1 \EXU/_2853_ ( .A(\_EXU_io_LSUIn_bits_wdata [9] ), .Z(\EXU/_0558_ ) );
BUF_X1 \EXU/_2854_ ( .A(\EXU/_0380_ ), .Z(\EXU/casez_tmp_0 [9] ) );
BUF_X1 \EXU/_2855_ ( .A(\EXU/in_imm [10] ), .Z(\EXU/_0396_ ) );
BUF_X1 \EXU/_2856_ ( .A(\_EXU_io_LSUIn_bits_wdata [10] ), .Z(\EXU/_0528_ ) );
BUF_X1 \EXU/_2857_ ( .A(\EXU/_0350_ ), .Z(\EXU/casez_tmp_0 [10] ) );
BUF_X1 \EXU/_2858_ ( .A(\EXU/in_imm [11] ), .Z(\EXU/_0397_ ) );
BUF_X1 \EXU/_2859_ ( .A(\_EXU_io_LSUIn_bits_wdata [11] ), .Z(\EXU/_0529_ ) );
BUF_X1 \EXU/_2860_ ( .A(\EXU/_0351_ ), .Z(\EXU/casez_tmp_0 [11] ) );
BUF_X1 \EXU/_2861_ ( .A(\EXU/in_imm [12] ), .Z(\EXU/_0398_ ) );
BUF_X1 \EXU/_2862_ ( .A(\_EXU_io_LSUIn_bits_wdata [12] ), .Z(\EXU/_0530_ ) );
BUF_X1 \EXU/_2863_ ( .A(\EXU/_0352_ ), .Z(\EXU/casez_tmp_0 [12] ) );
BUF_X1 \EXU/_2864_ ( .A(\EXU/in_imm [13] ), .Z(\EXU/_0399_ ) );
BUF_X1 \EXU/_2865_ ( .A(\_EXU_io_LSUIn_bits_wdata [13] ), .Z(\EXU/_0531_ ) );
BUF_X1 \EXU/_2866_ ( .A(\EXU/_0353_ ), .Z(\EXU/casez_tmp_0 [13] ) );
BUF_X1 \EXU/_2867_ ( .A(\EXU/in_imm [14] ), .Z(\EXU/_0400_ ) );
BUF_X1 \EXU/_2868_ ( .A(\_EXU_io_LSUIn_bits_wdata [14] ), .Z(\EXU/_0532_ ) );
BUF_X1 \EXU/_2869_ ( .A(\EXU/_0354_ ), .Z(\EXU/casez_tmp_0 [14] ) );
BUF_X1 \EXU/_2870_ ( .A(\EXU/in_imm [15] ), .Z(\EXU/_0401_ ) );
BUF_X1 \EXU/_2871_ ( .A(\_EXU_io_LSUIn_bits_wdata [15] ), .Z(\EXU/_0533_ ) );
BUF_X1 \EXU/_2872_ ( .A(\EXU/_0355_ ), .Z(\EXU/casez_tmp_0 [15] ) );
BUF_X1 \EXU/_2873_ ( .A(\EXU/in_imm [16] ), .Z(\EXU/_0402_ ) );
BUF_X1 \EXU/_2874_ ( .A(\_EXU_io_LSUIn_bits_wdata [16] ), .Z(\EXU/_0534_ ) );
BUF_X1 \EXU/_2875_ ( .A(\EXU/_0356_ ), .Z(\EXU/casez_tmp_0 [16] ) );
BUF_X1 \EXU/_2876_ ( .A(\EXU/in_imm [17] ), .Z(\EXU/_0403_ ) );
BUF_X1 \EXU/_2877_ ( .A(\_EXU_io_LSUIn_bits_wdata [17] ), .Z(\EXU/_0535_ ) );
BUF_X1 \EXU/_2878_ ( .A(\EXU/_0357_ ), .Z(\EXU/casez_tmp_0 [17] ) );
BUF_X1 \EXU/_2879_ ( .A(\EXU/in_imm [18] ), .Z(\EXU/_0404_ ) );
BUF_X1 \EXU/_2880_ ( .A(\_EXU_io_LSUIn_bits_wdata [18] ), .Z(\EXU/_0536_ ) );
BUF_X1 \EXU/_2881_ ( .A(\EXU/_0358_ ), .Z(\EXU/casez_tmp_0 [18] ) );
BUF_X1 \EXU/_2882_ ( .A(\EXU/in_imm [19] ), .Z(\EXU/_0405_ ) );
BUF_X1 \EXU/_2883_ ( .A(\_EXU_io_LSUIn_bits_wdata [19] ), .Z(\EXU/_0537_ ) );
BUF_X1 \EXU/_2884_ ( .A(\EXU/_0359_ ), .Z(\EXU/casez_tmp_0 [19] ) );
BUF_X1 \EXU/_2885_ ( .A(\EXU/in_imm [20] ), .Z(\EXU/_0407_ ) );
BUF_X1 \EXU/_2886_ ( .A(\_EXU_io_LSUIn_bits_wdata [20] ), .Z(\EXU/_0539_ ) );
BUF_X1 \EXU/_2887_ ( .A(\EXU/_0361_ ), .Z(\EXU/casez_tmp_0 [20] ) );
BUF_X1 \EXU/_2888_ ( .A(\EXU/in_imm [21] ), .Z(\EXU/_0408_ ) );
BUF_X1 \EXU/_2889_ ( .A(\_EXU_io_LSUIn_bits_wdata [21] ), .Z(\EXU/_0540_ ) );
BUF_X1 \EXU/_2890_ ( .A(\EXU/_0362_ ), .Z(\EXU/casez_tmp_0 [21] ) );
BUF_X1 \EXU/_2891_ ( .A(\EXU/in_imm [22] ), .Z(\EXU/_0409_ ) );
BUF_X1 \EXU/_2892_ ( .A(\_EXU_io_LSUIn_bits_wdata [22] ), .Z(\EXU/_0541_ ) );
BUF_X1 \EXU/_2893_ ( .A(\EXU/_0363_ ), .Z(\EXU/casez_tmp_0 [22] ) );
BUF_X1 \EXU/_2894_ ( .A(\EXU/in_imm [23] ), .Z(\EXU/_0410_ ) );
BUF_X1 \EXU/_2895_ ( .A(\_EXU_io_LSUIn_bits_wdata [23] ), .Z(\EXU/_0542_ ) );
BUF_X1 \EXU/_2896_ ( .A(\EXU/_0364_ ), .Z(\EXU/casez_tmp_0 [23] ) );
BUF_X1 \EXU/_2897_ ( .A(\EXU/in_imm [24] ), .Z(\EXU/_0411_ ) );
BUF_X1 \EXU/_2898_ ( .A(\_EXU_io_LSUIn_bits_wdata [24] ), .Z(\EXU/_0543_ ) );
BUF_X1 \EXU/_2899_ ( .A(\EXU/_0365_ ), .Z(\EXU/casez_tmp_0 [24] ) );
BUF_X1 \EXU/_2900_ ( .A(\EXU/in_imm [25] ), .Z(\EXU/_0412_ ) );
BUF_X1 \EXU/_2901_ ( .A(\_EXU_io_LSUIn_bits_wdata [25] ), .Z(\EXU/_0544_ ) );
BUF_X1 \EXU/_2902_ ( .A(\EXU/_0366_ ), .Z(\EXU/casez_tmp_0 [25] ) );
BUF_X1 \EXU/_2903_ ( .A(\EXU/in_imm [26] ), .Z(\EXU/_0413_ ) );
BUF_X1 \EXU/_2904_ ( .A(\_EXU_io_LSUIn_bits_wdata [26] ), .Z(\EXU/_0545_ ) );
BUF_X1 \EXU/_2905_ ( .A(\EXU/_0367_ ), .Z(\EXU/casez_tmp_0 [26] ) );
BUF_X1 \EXU/_2906_ ( .A(\EXU/in_imm [27] ), .Z(\EXU/_0414_ ) );
BUF_X1 \EXU/_2907_ ( .A(\_EXU_io_LSUIn_bits_wdata [27] ), .Z(\EXU/_0546_ ) );
BUF_X1 \EXU/_2908_ ( .A(\EXU/_0368_ ), .Z(\EXU/casez_tmp_0 [27] ) );
BUF_X1 \EXU/_2909_ ( .A(\EXU/in_imm [28] ), .Z(\EXU/_0415_ ) );
BUF_X1 \EXU/_2910_ ( .A(\_EXU_io_LSUIn_bits_wdata [28] ), .Z(\EXU/_0547_ ) );
BUF_X1 \EXU/_2911_ ( .A(\EXU/_0369_ ), .Z(\EXU/casez_tmp_0 [28] ) );
BUF_X1 \EXU/_2912_ ( .A(\EXU/in_imm [29] ), .Z(\EXU/_0416_ ) );
BUF_X1 \EXU/_2913_ ( .A(\_EXU_io_LSUIn_bits_wdata [29] ), .Z(\EXU/_0548_ ) );
BUF_X1 \EXU/_2914_ ( .A(\EXU/_0370_ ), .Z(\EXU/casez_tmp_0 [29] ) );
BUF_X1 \EXU/_2915_ ( .A(\EXU/in_imm [30] ), .Z(\EXU/_0418_ ) );
BUF_X1 \EXU/_2916_ ( .A(\_EXU_io_LSUIn_bits_wdata [30] ), .Z(\EXU/_0550_ ) );
BUF_X1 \EXU/_2917_ ( .A(\EXU/_0372_ ), .Z(\EXU/casez_tmp_0 [30] ) );
BUF_X1 \EXU/_2918_ ( .A(\EXU/in_imm [31] ), .Z(\EXU/_0419_ ) );
BUF_X1 \EXU/_2919_ ( .A(\_EXU_io_LSUIn_bits_wdata [31] ), .Z(\EXU/_0551_ ) );
BUF_X1 \EXU/_2920_ ( .A(\EXU/_0373_ ), .Z(\EXU/casez_tmp_0 [31] ) );
BUF_X1 \EXU/_2921_ ( .A(_WBU_io_in_ready ), .Z(\EXU/_0841_ ) );
BUF_X1 \EXU/_2922_ ( .A(_LSU_io_out_valid ), .Z(\EXU/_0595_ ) );
BUF_X1 \EXU/_2923_ ( .A(_LSU_io_in_ready ), .Z(\EXU/_0560_ ) );
BUF_X1 \EXU/_2924_ ( .A(_IDU_io_out_bits_control_memRen ), .Z(\EXU/_0613_ ) );
BUF_X1 \EXU/_2925_ ( .A(_IDU_io_out_bits_control_memWen ), .Z(\EXU/_0614_ ) );
BUF_X1 \EXU/_2926_ ( .A(\EXU/_BrCond_io_PCASrc ), .Z(\EXU/_0067_ ) );
BUF_X1 \EXU/_2927_ ( .A(\EXU/_BrCond_io_PCBSrc ), .Z(\EXU/_0068_ ) );
BUF_X1 \EXU/_2928_ ( .A(\EXU/_0820_ ), .Z(\_EXU_io_out_bits_pcCom [1] ) );
BUF_X1 \EXU/_2929_ ( .A(\EXU/_0831_ ), .Z(\_EXU_io_out_bits_pcCom [2] ) );
BUF_X1 \EXU/_2930_ ( .A(\EXU/_0834_ ), .Z(\_EXU_io_out_bits_pcCom [3] ) );
BUF_X1 \EXU/_2931_ ( .A(\EXU/_0835_ ), .Z(\_EXU_io_out_bits_pcCom [4] ) );
BUF_X1 \EXU/_2932_ ( .A(\EXU/_0836_ ), .Z(\_EXU_io_out_bits_pcCom [5] ) );
BUF_X1 \EXU/_2933_ ( .A(\EXU/_0837_ ), .Z(\_EXU_io_out_bits_pcCom [6] ) );
BUF_X1 \EXU/_2934_ ( .A(\EXU/_0838_ ), .Z(\_EXU_io_out_bits_pcCom [7] ) );
BUF_X1 \EXU/_2935_ ( .A(\EXU/_0839_ ), .Z(\_EXU_io_out_bits_pcCom [8] ) );
BUF_X1 \EXU/_2936_ ( .A(\EXU/_0840_ ), .Z(\_EXU_io_out_bits_pcCom [9] ) );
BUF_X1 \EXU/_2937_ ( .A(\EXU/_0810_ ), .Z(\_EXU_io_out_bits_pcCom [10] ) );
BUF_X1 \EXU/_2938_ ( .A(\EXU/_0811_ ), .Z(\_EXU_io_out_bits_pcCom [11] ) );
BUF_X1 \EXU/_2939_ ( .A(\EXU/_0812_ ), .Z(\_EXU_io_out_bits_pcCom [12] ) );
BUF_X1 \EXU/_2940_ ( .A(\EXU/_0813_ ), .Z(\_EXU_io_out_bits_pcCom [13] ) );
BUF_X1 \EXU/_2941_ ( .A(\EXU/_0814_ ), .Z(\_EXU_io_out_bits_pcCom [14] ) );
BUF_X1 \EXU/_2942_ ( .A(\EXU/_0815_ ), .Z(\_EXU_io_out_bits_pcCom [15] ) );
BUF_X1 \EXU/_2943_ ( .A(\EXU/_0816_ ), .Z(\_EXU_io_out_bits_pcCom [16] ) );
BUF_X1 \EXU/_2944_ ( .A(\EXU/_0817_ ), .Z(\_EXU_io_out_bits_pcCom [17] ) );
BUF_X1 \EXU/_2945_ ( .A(\EXU/_0818_ ), .Z(\_EXU_io_out_bits_pcCom [18] ) );
BUF_X1 \EXU/_2946_ ( .A(\EXU/_0819_ ), .Z(\_EXU_io_out_bits_pcCom [19] ) );
BUF_X1 \EXU/_2947_ ( .A(\EXU/_0821_ ), .Z(\_EXU_io_out_bits_pcCom [20] ) );
BUF_X1 \EXU/_2948_ ( .A(\EXU/_0822_ ), .Z(\_EXU_io_out_bits_pcCom [21] ) );
BUF_X1 \EXU/_2949_ ( .A(\EXU/_0823_ ), .Z(\_EXU_io_out_bits_pcCom [22] ) );
BUF_X1 \EXU/_2950_ ( .A(\EXU/_0824_ ), .Z(\_EXU_io_out_bits_pcCom [23] ) );
BUF_X1 \EXU/_2951_ ( .A(\EXU/_0825_ ), .Z(\_EXU_io_out_bits_pcCom [24] ) );
BUF_X1 \EXU/_2952_ ( .A(\EXU/_0826_ ), .Z(\_EXU_io_out_bits_pcCom [25] ) );
BUF_X1 \EXU/_2953_ ( .A(\EXU/_0827_ ), .Z(\_EXU_io_out_bits_pcCom [26] ) );
BUF_X1 \EXU/_2954_ ( .A(\EXU/_0828_ ), .Z(\_EXU_io_out_bits_pcCom [27] ) );
BUF_X1 \EXU/_2955_ ( .A(\EXU/_0829_ ), .Z(\_EXU_io_out_bits_pcCom [28] ) );
BUF_X1 \EXU/_2956_ ( .A(\EXU/_0830_ ), .Z(\_EXU_io_out_bits_pcCom [29] ) );
BUF_X1 \EXU/_2957_ ( .A(\EXU/_0832_ ), .Z(\_EXU_io_out_bits_pcCom [30] ) );
BUF_X1 \EXU/_2958_ ( .A(\EXU/_0833_ ), .Z(\_EXU_io_out_bits_pcCom [31] ) );
BUF_X1 \EXU/_2959_ ( .A(\EXU/_0809_ ), .Z(\_EXU_io_out_bits_pcCom [0] ) );
BUF_X1 \EXU/_2960_ ( .A(\_EXU_io_out_bits_memOut [0] ), .Z(\EXU/_0777_ ) );
BUF_X1 \EXU/_2961_ ( .A(\_LSU_io_out_bits_rdata [0] ), .Z(\EXU/_0562_ ) );
BUF_X1 \EXU/_2962_ ( .A(\EXU/_0136_ ), .Z(\EXU/_1430_ ) );
BUF_X1 \EXU/_2963_ ( .A(\_EXU_io_out_bits_memOut [1] ), .Z(\EXU/_0788_ ) );
BUF_X1 \EXU/_2964_ ( .A(\_LSU_io_out_bits_rdata [1] ), .Z(\EXU/_0573_ ) );
BUF_X1 \EXU/_2965_ ( .A(\EXU/_0137_ ), .Z(\EXU/_1431_ ) );
BUF_X1 \EXU/_2966_ ( .A(\_EXU_io_out_bits_memOut [2] ), .Z(\EXU/_0799_ ) );
BUF_X1 \EXU/_2967_ ( .A(\_LSU_io_out_bits_rdata [2] ), .Z(\EXU/_0584_ ) );
BUF_X1 \EXU/_2968_ ( .A(\EXU/_0138_ ), .Z(\EXU/_1432_ ) );
BUF_X1 \EXU/_2969_ ( .A(\_EXU_io_out_bits_memOut [3] ), .Z(\EXU/_0802_ ) );
BUF_X1 \EXU/_2970_ ( .A(\_LSU_io_out_bits_rdata [3] ), .Z(\EXU/_0587_ ) );
BUF_X1 \EXU/_2971_ ( .A(\EXU/_0139_ ), .Z(\EXU/_1433_ ) );
BUF_X1 \EXU/_2972_ ( .A(\_EXU_io_out_bits_memOut [4] ), .Z(\EXU/_0803_ ) );
BUF_X1 \EXU/_2973_ ( .A(\_LSU_io_out_bits_rdata [4] ), .Z(\EXU/_0588_ ) );
BUF_X1 \EXU/_2974_ ( .A(\EXU/_0140_ ), .Z(\EXU/_1434_ ) );
BUF_X1 \EXU/_2975_ ( .A(\_EXU_io_out_bits_memOut [5] ), .Z(\EXU/_0804_ ) );
BUF_X1 \EXU/_2976_ ( .A(\_LSU_io_out_bits_rdata [5] ), .Z(\EXU/_0589_ ) );
BUF_X1 \EXU/_2977_ ( .A(\EXU/_0141_ ), .Z(\EXU/_1435_ ) );
BUF_X1 \EXU/_2978_ ( .A(\_EXU_io_out_bits_memOut [6] ), .Z(\EXU/_0805_ ) );
BUF_X1 \EXU/_2979_ ( .A(\_LSU_io_out_bits_rdata [6] ), .Z(\EXU/_0590_ ) );
BUF_X1 \EXU/_2980_ ( .A(\EXU/_0142_ ), .Z(\EXU/_1436_ ) );
BUF_X1 \EXU/_2981_ ( .A(\_EXU_io_out_bits_memOut [7] ), .Z(\EXU/_0806_ ) );
BUF_X1 \EXU/_2982_ ( .A(\_LSU_io_out_bits_rdata [7] ), .Z(\EXU/_0591_ ) );
BUF_X1 \EXU/_2983_ ( .A(\EXU/_0143_ ), .Z(\EXU/_1437_ ) );
BUF_X1 \EXU/_2984_ ( .A(\_EXU_io_out_bits_memOut [8] ), .Z(\EXU/_0807_ ) );
BUF_X1 \EXU/_2985_ ( .A(\_LSU_io_out_bits_rdata [8] ), .Z(\EXU/_0592_ ) );
BUF_X1 \EXU/_2986_ ( .A(\EXU/_0144_ ), .Z(\EXU/_1438_ ) );
BUF_X1 \EXU/_2987_ ( .A(\_EXU_io_out_bits_memOut [9] ), .Z(\EXU/_0808_ ) );
BUF_X1 \EXU/_2988_ ( .A(\_LSU_io_out_bits_rdata [9] ), .Z(\EXU/_0593_ ) );
BUF_X1 \EXU/_2989_ ( .A(\EXU/_0145_ ), .Z(\EXU/_1439_ ) );
BUF_X1 \EXU/_2990_ ( .A(\_EXU_io_out_bits_memOut [10] ), .Z(\EXU/_0778_ ) );
BUF_X1 \EXU/_2991_ ( .A(\_LSU_io_out_bits_rdata [10] ), .Z(\EXU/_0563_ ) );
BUF_X1 \EXU/_2992_ ( .A(\EXU/_0146_ ), .Z(\EXU/_1440_ ) );
BUF_X1 \EXU/_2993_ ( .A(\_EXU_io_out_bits_memOut [11] ), .Z(\EXU/_0779_ ) );
BUF_X1 \EXU/_2994_ ( .A(\_LSU_io_out_bits_rdata [11] ), .Z(\EXU/_0564_ ) );
BUF_X1 \EXU/_2995_ ( .A(\EXU/_0147_ ), .Z(\EXU/_1441_ ) );
BUF_X1 \EXU/_2996_ ( .A(\_EXU_io_out_bits_memOut [12] ), .Z(\EXU/_0780_ ) );
BUF_X1 \EXU/_2997_ ( .A(\_LSU_io_out_bits_rdata [12] ), .Z(\EXU/_0565_ ) );
BUF_X1 \EXU/_2998_ ( .A(\EXU/_0148_ ), .Z(\EXU/_1442_ ) );
BUF_X1 \EXU/_2999_ ( .A(\_EXU_io_out_bits_memOut [13] ), .Z(\EXU/_0781_ ) );
BUF_X1 \EXU/_3000_ ( .A(\_LSU_io_out_bits_rdata [13] ), .Z(\EXU/_0566_ ) );
BUF_X1 \EXU/_3001_ ( .A(\EXU/_0149_ ), .Z(\EXU/_1443_ ) );
BUF_X1 \EXU/_3002_ ( .A(\_EXU_io_out_bits_memOut [14] ), .Z(\EXU/_0782_ ) );
BUF_X1 \EXU/_3003_ ( .A(\_LSU_io_out_bits_rdata [14] ), .Z(\EXU/_0567_ ) );
BUF_X1 \EXU/_3004_ ( .A(\EXU/_0150_ ), .Z(\EXU/_1444_ ) );
BUF_X1 \EXU/_3005_ ( .A(\_EXU_io_out_bits_memOut [15] ), .Z(\EXU/_0783_ ) );
BUF_X1 \EXU/_3006_ ( .A(\_LSU_io_out_bits_rdata [15] ), .Z(\EXU/_0568_ ) );
BUF_X1 \EXU/_3007_ ( .A(\EXU/_0151_ ), .Z(\EXU/_1445_ ) );
BUF_X1 \EXU/_3008_ ( .A(\_EXU_io_out_bits_memOut [16] ), .Z(\EXU/_0784_ ) );
BUF_X1 \EXU/_3009_ ( .A(\_LSU_io_out_bits_rdata [16] ), .Z(\EXU/_0569_ ) );
BUF_X1 \EXU/_3010_ ( .A(\EXU/_0152_ ), .Z(\EXU/_1446_ ) );
BUF_X1 \EXU/_3011_ ( .A(\_EXU_io_out_bits_memOut [17] ), .Z(\EXU/_0785_ ) );
BUF_X1 \EXU/_3012_ ( .A(\_LSU_io_out_bits_rdata [17] ), .Z(\EXU/_0570_ ) );
BUF_X1 \EXU/_3013_ ( .A(\EXU/_0153_ ), .Z(\EXU/_1447_ ) );
BUF_X1 \EXU/_3014_ ( .A(\_EXU_io_out_bits_memOut [18] ), .Z(\EXU/_0786_ ) );
BUF_X1 \EXU/_3015_ ( .A(\_LSU_io_out_bits_rdata [18] ), .Z(\EXU/_0571_ ) );
BUF_X1 \EXU/_3016_ ( .A(\EXU/_0154_ ), .Z(\EXU/_1448_ ) );
BUF_X1 \EXU/_3017_ ( .A(\_EXU_io_out_bits_memOut [19] ), .Z(\EXU/_0787_ ) );
BUF_X1 \EXU/_3018_ ( .A(\_LSU_io_out_bits_rdata [19] ), .Z(\EXU/_0572_ ) );
BUF_X1 \EXU/_3019_ ( .A(\EXU/_0155_ ), .Z(\EXU/_1449_ ) );
BUF_X1 \EXU/_3020_ ( .A(\_EXU_io_out_bits_memOut [20] ), .Z(\EXU/_0789_ ) );
BUF_X1 \EXU/_3021_ ( .A(\_LSU_io_out_bits_rdata [20] ), .Z(\EXU/_0574_ ) );
BUF_X1 \EXU/_3022_ ( .A(\EXU/_0156_ ), .Z(\EXU/_1450_ ) );
BUF_X1 \EXU/_3023_ ( .A(\_EXU_io_out_bits_memOut [21] ), .Z(\EXU/_0790_ ) );
BUF_X1 \EXU/_3024_ ( .A(\_LSU_io_out_bits_rdata [21] ), .Z(\EXU/_0575_ ) );
BUF_X1 \EXU/_3025_ ( .A(\EXU/_0157_ ), .Z(\EXU/_1451_ ) );
BUF_X1 \EXU/_3026_ ( .A(\_EXU_io_out_bits_memOut [22] ), .Z(\EXU/_0791_ ) );
BUF_X1 \EXU/_3027_ ( .A(\_LSU_io_out_bits_rdata [22] ), .Z(\EXU/_0576_ ) );
BUF_X1 \EXU/_3028_ ( .A(\EXU/_0158_ ), .Z(\EXU/_1452_ ) );
BUF_X1 \EXU/_3029_ ( .A(\_EXU_io_out_bits_memOut [23] ), .Z(\EXU/_0792_ ) );
BUF_X1 \EXU/_3030_ ( .A(\_LSU_io_out_bits_rdata [23] ), .Z(\EXU/_0577_ ) );
BUF_X1 \EXU/_3031_ ( .A(\EXU/_0159_ ), .Z(\EXU/_1453_ ) );
BUF_X1 \EXU/_3032_ ( .A(\_EXU_io_out_bits_memOut [24] ), .Z(\EXU/_0793_ ) );
BUF_X1 \EXU/_3033_ ( .A(\_LSU_io_out_bits_rdata [24] ), .Z(\EXU/_0578_ ) );
BUF_X1 \EXU/_3034_ ( .A(\EXU/_0160_ ), .Z(\EXU/_1454_ ) );
BUF_X1 \EXU/_3035_ ( .A(\_EXU_io_out_bits_memOut [25] ), .Z(\EXU/_0794_ ) );
BUF_X1 \EXU/_3036_ ( .A(\_LSU_io_out_bits_rdata [25] ), .Z(\EXU/_0579_ ) );
BUF_X1 \EXU/_3037_ ( .A(\EXU/_0161_ ), .Z(\EXU/_1455_ ) );
BUF_X1 \EXU/_3038_ ( .A(\_EXU_io_out_bits_memOut [26] ), .Z(\EXU/_0795_ ) );
BUF_X1 \EXU/_3039_ ( .A(\_LSU_io_out_bits_rdata [26] ), .Z(\EXU/_0580_ ) );
BUF_X1 \EXU/_3040_ ( .A(\EXU/_0162_ ), .Z(\EXU/_1456_ ) );
BUF_X1 \EXU/_3041_ ( .A(\_EXU_io_out_bits_memOut [27] ), .Z(\EXU/_0796_ ) );
BUF_X1 \EXU/_3042_ ( .A(\_LSU_io_out_bits_rdata [27] ), .Z(\EXU/_0581_ ) );
BUF_X1 \EXU/_3043_ ( .A(\EXU/_0163_ ), .Z(\EXU/_1457_ ) );
BUF_X1 \EXU/_3044_ ( .A(\_EXU_io_out_bits_memOut [28] ), .Z(\EXU/_0797_ ) );
BUF_X1 \EXU/_3045_ ( .A(\_LSU_io_out_bits_rdata [28] ), .Z(\EXU/_0582_ ) );
BUF_X1 \EXU/_3046_ ( .A(\EXU/_0164_ ), .Z(\EXU/_1458_ ) );
BUF_X1 \EXU/_3047_ ( .A(\_EXU_io_out_bits_memOut [29] ), .Z(\EXU/_0798_ ) );
BUF_X1 \EXU/_3048_ ( .A(\_LSU_io_out_bits_rdata [29] ), .Z(\EXU/_0583_ ) );
BUF_X1 \EXU/_3049_ ( .A(\EXU/_0165_ ), .Z(\EXU/_1459_ ) );
BUF_X1 \EXU/_3050_ ( .A(\_EXU_io_out_bits_memOut [30] ), .Z(\EXU/_0800_ ) );
BUF_X1 \EXU/_3051_ ( .A(\_LSU_io_out_bits_rdata [30] ), .Z(\EXU/_0585_ ) );
BUF_X1 \EXU/_3052_ ( .A(\EXU/_0166_ ), .Z(\EXU/_1460_ ) );
BUF_X1 \EXU/_3053_ ( .A(\_EXU_io_out_bits_memOut [31] ), .Z(\EXU/_0801_ ) );
BUF_X1 \EXU/_3054_ ( .A(\_LSU_io_out_bits_rdata [31] ), .Z(\EXU/_0586_ ) );
BUF_X1 \EXU/_3055_ ( .A(\EXU/_0167_ ), .Z(\EXU/_1461_ ) );
BUF_X1 \EXU/_3056_ ( .A(\_IDU_io_out_bits_pc [0] ), .Z(\EXU/_0647_ ) );
BUF_X1 \EXU/_3057_ ( .A(\EXU/_0170_ ), .Z(\EXU/_1464_ ) );
BUF_X1 \EXU/_3058_ ( .A(\_IDU_io_out_bits_pc [1] ), .Z(\EXU/_0658_ ) );
BUF_X1 \EXU/_3059_ ( .A(\EXU/_0171_ ), .Z(\EXU/_1465_ ) );
BUF_X1 \EXU/_3060_ ( .A(\_IDU_io_out_bits_pc [2] ), .Z(\EXU/_0669_ ) );
BUF_X1 \EXU/_3061_ ( .A(\EXU/_0172_ ), .Z(\EXU/_1466_ ) );
BUF_X1 \EXU/_3062_ ( .A(\_IDU_io_out_bits_pc [3] ), .Z(\EXU/_0672_ ) );
BUF_X1 \EXU/_3063_ ( .A(\EXU/_0173_ ), .Z(\EXU/_1467_ ) );
BUF_X1 \EXU/_3064_ ( .A(\_IDU_io_out_bits_pc [4] ), .Z(\EXU/_0673_ ) );
BUF_X1 \EXU/_3065_ ( .A(\EXU/_0174_ ), .Z(\EXU/_1468_ ) );
BUF_X1 \EXU/_3066_ ( .A(\_IDU_io_out_bits_pc [5] ), .Z(\EXU/_0674_ ) );
BUF_X1 \EXU/_3067_ ( .A(\EXU/_0175_ ), .Z(\EXU/_1469_ ) );
BUF_X1 \EXU/_3068_ ( .A(\_IDU_io_out_bits_pc [6] ), .Z(\EXU/_0675_ ) );
BUF_X1 \EXU/_3069_ ( .A(\EXU/_0176_ ), .Z(\EXU/_1470_ ) );
BUF_X1 \EXU/_3070_ ( .A(\_IDU_io_out_bits_pc [7] ), .Z(\EXU/_0676_ ) );
BUF_X1 \EXU/_3071_ ( .A(\EXU/_0177_ ), .Z(\EXU/_1471_ ) );
BUF_X1 \EXU/_3072_ ( .A(\_IDU_io_out_bits_pc [8] ), .Z(\EXU/_0677_ ) );
BUF_X1 \EXU/_3073_ ( .A(\EXU/_0178_ ), .Z(\EXU/_1472_ ) );
BUF_X1 \EXU/_3074_ ( .A(\_IDU_io_out_bits_pc [9] ), .Z(\EXU/_0678_ ) );
BUF_X1 \EXU/_3075_ ( .A(\EXU/_0179_ ), .Z(\EXU/_1473_ ) );
BUF_X1 \EXU/_3076_ ( .A(\_IDU_io_out_bits_pc [10] ), .Z(\EXU/_0648_ ) );
BUF_X1 \EXU/_3077_ ( .A(\EXU/_0180_ ), .Z(\EXU/_1474_ ) );
BUF_X1 \EXU/_3078_ ( .A(\_IDU_io_out_bits_pc [11] ), .Z(\EXU/_0649_ ) );
BUF_X1 \EXU/_3079_ ( .A(\EXU/_0181_ ), .Z(\EXU/_1475_ ) );
BUF_X1 \EXU/_3080_ ( .A(\_IDU_io_out_bits_pc [12] ), .Z(\EXU/_0650_ ) );
BUF_X1 \EXU/_3081_ ( .A(\EXU/_0182_ ), .Z(\EXU/_1476_ ) );
BUF_X1 \EXU/_3082_ ( .A(\_IDU_io_out_bits_pc [13] ), .Z(\EXU/_0651_ ) );
BUF_X1 \EXU/_3083_ ( .A(\EXU/_0183_ ), .Z(\EXU/_1477_ ) );
BUF_X1 \EXU/_3084_ ( .A(\_IDU_io_out_bits_pc [14] ), .Z(\EXU/_0652_ ) );
BUF_X1 \EXU/_3085_ ( .A(\EXU/_0184_ ), .Z(\EXU/_1478_ ) );
BUF_X1 \EXU/_3086_ ( .A(\_IDU_io_out_bits_pc [15] ), .Z(\EXU/_0653_ ) );
BUF_X1 \EXU/_3087_ ( .A(\EXU/_0185_ ), .Z(\EXU/_1479_ ) );
BUF_X1 \EXU/_3088_ ( .A(\_IDU_io_out_bits_pc [16] ), .Z(\EXU/_0654_ ) );
BUF_X1 \EXU/_3089_ ( .A(\EXU/_0186_ ), .Z(\EXU/_1480_ ) );
BUF_X1 \EXU/_3090_ ( .A(\_IDU_io_out_bits_pc [17] ), .Z(\EXU/_0655_ ) );
BUF_X1 \EXU/_3091_ ( .A(\EXU/_0187_ ), .Z(\EXU/_1481_ ) );
BUF_X1 \EXU/_3092_ ( .A(\_IDU_io_out_bits_pc [18] ), .Z(\EXU/_0656_ ) );
BUF_X1 \EXU/_3093_ ( .A(\EXU/_0188_ ), .Z(\EXU/_1482_ ) );
BUF_X1 \EXU/_3094_ ( .A(\_IDU_io_out_bits_pc [19] ), .Z(\EXU/_0657_ ) );
BUF_X1 \EXU/_3095_ ( .A(\EXU/_0189_ ), .Z(\EXU/_1483_ ) );
BUF_X1 \EXU/_3096_ ( .A(\_IDU_io_out_bits_pc [20] ), .Z(\EXU/_0659_ ) );
BUF_X1 \EXU/_3097_ ( .A(\EXU/_0190_ ), .Z(\EXU/_1484_ ) );
BUF_X1 \EXU/_3098_ ( .A(\_IDU_io_out_bits_pc [21] ), .Z(\EXU/_0660_ ) );
BUF_X1 \EXU/_3099_ ( .A(\EXU/_0191_ ), .Z(\EXU/_1485_ ) );
BUF_X1 \EXU/_3100_ ( .A(\_IDU_io_out_bits_pc [22] ), .Z(\EXU/_0661_ ) );
BUF_X1 \EXU/_3101_ ( .A(\EXU/_0192_ ), .Z(\EXU/_1486_ ) );
BUF_X1 \EXU/_3102_ ( .A(\_IDU_io_out_bits_pc [23] ), .Z(\EXU/_0662_ ) );
BUF_X1 \EXU/_3103_ ( .A(\EXU/_0193_ ), .Z(\EXU/_1487_ ) );
BUF_X1 \EXU/_3104_ ( .A(\_IDU_io_out_bits_pc [24] ), .Z(\EXU/_0663_ ) );
BUF_X1 \EXU/_3105_ ( .A(\EXU/_0194_ ), .Z(\EXU/_1488_ ) );
BUF_X1 \EXU/_3106_ ( .A(\_IDU_io_out_bits_pc [25] ), .Z(\EXU/_0664_ ) );
BUF_X1 \EXU/_3107_ ( .A(\EXU/_0195_ ), .Z(\EXU/_1489_ ) );
BUF_X1 \EXU/_3108_ ( .A(\_IDU_io_out_bits_pc [26] ), .Z(\EXU/_0665_ ) );
BUF_X1 \EXU/_3109_ ( .A(\EXU/_0196_ ), .Z(\EXU/_1490_ ) );
BUF_X1 \EXU/_3110_ ( .A(\_IDU_io_out_bits_pc [27] ), .Z(\EXU/_0666_ ) );
BUF_X1 \EXU/_3111_ ( .A(\EXU/_0197_ ), .Z(\EXU/_1491_ ) );
BUF_X1 \EXU/_3112_ ( .A(\_IDU_io_out_bits_pc [28] ), .Z(\EXU/_0667_ ) );
BUF_X1 \EXU/_3113_ ( .A(\EXU/_0198_ ), .Z(\EXU/_1492_ ) );
BUF_X1 \EXU/_3114_ ( .A(\_IDU_io_out_bits_pc [29] ), .Z(\EXU/_0668_ ) );
BUF_X1 \EXU/_3115_ ( .A(\EXU/_0199_ ), .Z(\EXU/_1493_ ) );
BUF_X1 \EXU/_3116_ ( .A(\_IDU_io_out_bits_pc [30] ), .Z(\EXU/_0670_ ) );
BUF_X1 \EXU/_3117_ ( .A(\EXU/_0200_ ), .Z(\EXU/_1494_ ) );
BUF_X1 \EXU/_3118_ ( .A(\_IDU_io_out_bits_pc [31] ), .Z(\EXU/_0671_ ) );
BUF_X1 \EXU/_3119_ ( .A(\EXU/_0201_ ), .Z(\EXU/_1495_ ) );
BUF_X1 \EXU/_3120_ ( .A(\_IDU_io_out_bits_rd1 [0] ), .Z(\EXU/_0679_ ) );
BUF_X1 \EXU/_3121_ ( .A(\EXU/_0202_ ), .Z(\EXU/_1496_ ) );
BUF_X1 \EXU/_3122_ ( .A(\_IDU_io_out_bits_rd1 [1] ), .Z(\EXU/_0690_ ) );
BUF_X1 \EXU/_3123_ ( .A(\EXU/_0203_ ), .Z(\EXU/_1497_ ) );
BUF_X1 \EXU/_3124_ ( .A(\_IDU_io_out_bits_rd1 [2] ), .Z(\EXU/_0701_ ) );
BUF_X1 \EXU/_3125_ ( .A(\EXU/_0204_ ), .Z(\EXU/_1498_ ) );
BUF_X1 \EXU/_3126_ ( .A(\_IDU_io_out_bits_rd1 [3] ), .Z(\EXU/_0704_ ) );
BUF_X1 \EXU/_3127_ ( .A(\EXU/_0205_ ), .Z(\EXU/_1499_ ) );
BUF_X1 \EXU/_3128_ ( .A(\_IDU_io_out_bits_rd1 [4] ), .Z(\EXU/_0705_ ) );
BUF_X1 \EXU/_3129_ ( .A(\EXU/_0206_ ), .Z(\EXU/_1500_ ) );
BUF_X1 \EXU/_3130_ ( .A(\_IDU_io_out_bits_rd1 [5] ), .Z(\EXU/_0706_ ) );
BUF_X1 \EXU/_3131_ ( .A(\EXU/_0207_ ), .Z(\EXU/_1501_ ) );
BUF_X1 \EXU/_3132_ ( .A(\_IDU_io_out_bits_rd1 [6] ), .Z(\EXU/_0707_ ) );
BUF_X1 \EXU/_3133_ ( .A(\EXU/_0208_ ), .Z(\EXU/_1502_ ) );
BUF_X1 \EXU/_3134_ ( .A(\_IDU_io_out_bits_rd1 [7] ), .Z(\EXU/_0708_ ) );
BUF_X1 \EXU/_3135_ ( .A(\EXU/_0209_ ), .Z(\EXU/_1503_ ) );
BUF_X1 \EXU/_3136_ ( .A(\_IDU_io_out_bits_rd1 [8] ), .Z(\EXU/_0709_ ) );
BUF_X1 \EXU/_3137_ ( .A(\EXU/_0210_ ), .Z(\EXU/_1504_ ) );
BUF_X1 \EXU/_3138_ ( .A(\_IDU_io_out_bits_rd1 [9] ), .Z(\EXU/_0710_ ) );
BUF_X1 \EXU/_3139_ ( .A(\EXU/_0211_ ), .Z(\EXU/_1505_ ) );
BUF_X1 \EXU/_3140_ ( .A(\_IDU_io_out_bits_rd1 [10] ), .Z(\EXU/_0680_ ) );
BUF_X1 \EXU/_3141_ ( .A(\EXU/_0212_ ), .Z(\EXU/_1506_ ) );
BUF_X1 \EXU/_3142_ ( .A(\_IDU_io_out_bits_rd1 [11] ), .Z(\EXU/_0681_ ) );
BUF_X1 \EXU/_3143_ ( .A(\EXU/_0213_ ), .Z(\EXU/_1507_ ) );
BUF_X1 \EXU/_3144_ ( .A(\_IDU_io_out_bits_rd1 [12] ), .Z(\EXU/_0682_ ) );
BUF_X1 \EXU/_3145_ ( .A(\EXU/_0214_ ), .Z(\EXU/_1508_ ) );
BUF_X1 \EXU/_3146_ ( .A(\_IDU_io_out_bits_rd1 [13] ), .Z(\EXU/_0683_ ) );
BUF_X1 \EXU/_3147_ ( .A(\EXU/_0215_ ), .Z(\EXU/_1509_ ) );
BUF_X1 \EXU/_3148_ ( .A(\_IDU_io_out_bits_rd1 [14] ), .Z(\EXU/_0684_ ) );
BUF_X1 \EXU/_3149_ ( .A(\EXU/_0216_ ), .Z(\EXU/_1510_ ) );
BUF_X1 \EXU/_3150_ ( .A(\_IDU_io_out_bits_rd1 [15] ), .Z(\EXU/_0685_ ) );
BUF_X1 \EXU/_3151_ ( .A(\EXU/_0217_ ), .Z(\EXU/_1511_ ) );
BUF_X1 \EXU/_3152_ ( .A(\_IDU_io_out_bits_rd1 [16] ), .Z(\EXU/_0686_ ) );
BUF_X1 \EXU/_3153_ ( .A(\EXU/_0218_ ), .Z(\EXU/_1512_ ) );
BUF_X1 \EXU/_3154_ ( .A(\_IDU_io_out_bits_rd1 [17] ), .Z(\EXU/_0687_ ) );
BUF_X1 \EXU/_3155_ ( .A(\EXU/_0219_ ), .Z(\EXU/_1513_ ) );
BUF_X1 \EXU/_3156_ ( .A(\_IDU_io_out_bits_rd1 [18] ), .Z(\EXU/_0688_ ) );
BUF_X1 \EXU/_3157_ ( .A(\EXU/_0220_ ), .Z(\EXU/_1514_ ) );
BUF_X1 \EXU/_3158_ ( .A(\_IDU_io_out_bits_rd1 [19] ), .Z(\EXU/_0689_ ) );
BUF_X1 \EXU/_3159_ ( .A(\EXU/_0221_ ), .Z(\EXU/_1515_ ) );
BUF_X1 \EXU/_3160_ ( .A(\_IDU_io_out_bits_rd1 [20] ), .Z(\EXU/_0691_ ) );
BUF_X1 \EXU/_3161_ ( .A(\EXU/_0222_ ), .Z(\EXU/_1516_ ) );
BUF_X1 \EXU/_3162_ ( .A(\_IDU_io_out_bits_rd1 [21] ), .Z(\EXU/_0692_ ) );
BUF_X1 \EXU/_3163_ ( .A(\EXU/_0223_ ), .Z(\EXU/_1517_ ) );
BUF_X1 \EXU/_3164_ ( .A(\_IDU_io_out_bits_rd1 [22] ), .Z(\EXU/_0693_ ) );
BUF_X1 \EXU/_3165_ ( .A(\EXU/_0224_ ), .Z(\EXU/_1518_ ) );
BUF_X1 \EXU/_3166_ ( .A(\_IDU_io_out_bits_rd1 [23] ), .Z(\EXU/_0694_ ) );
BUF_X1 \EXU/_3167_ ( .A(\EXU/_0225_ ), .Z(\EXU/_1519_ ) );
BUF_X1 \EXU/_3168_ ( .A(\_IDU_io_out_bits_rd1 [24] ), .Z(\EXU/_0695_ ) );
BUF_X1 \EXU/_3169_ ( .A(\EXU/_0226_ ), .Z(\EXU/_1520_ ) );
BUF_X1 \EXU/_3170_ ( .A(\_IDU_io_out_bits_rd1 [25] ), .Z(\EXU/_0696_ ) );
BUF_X1 \EXU/_3171_ ( .A(\EXU/_0227_ ), .Z(\EXU/_1521_ ) );
BUF_X1 \EXU/_3172_ ( .A(\_IDU_io_out_bits_rd1 [26] ), .Z(\EXU/_0697_ ) );
BUF_X1 \EXU/_3173_ ( .A(\EXU/_0228_ ), .Z(\EXU/_1522_ ) );
BUF_X1 \EXU/_3174_ ( .A(\_IDU_io_out_bits_rd1 [27] ), .Z(\EXU/_0698_ ) );
BUF_X1 \EXU/_3175_ ( .A(\EXU/_0229_ ), .Z(\EXU/_1523_ ) );
BUF_X1 \EXU/_3176_ ( .A(\_IDU_io_out_bits_rd1 [28] ), .Z(\EXU/_0699_ ) );
BUF_X1 \EXU/_3177_ ( .A(\EXU/_0230_ ), .Z(\EXU/_1524_ ) );
BUF_X1 \EXU/_3178_ ( .A(\_IDU_io_out_bits_rd1 [29] ), .Z(\EXU/_0700_ ) );
BUF_X1 \EXU/_3179_ ( .A(\EXU/_0231_ ), .Z(\EXU/_1525_ ) );
BUF_X1 \EXU/_3180_ ( .A(\_IDU_io_out_bits_rd1 [30] ), .Z(\EXU/_0702_ ) );
BUF_X1 \EXU/_3181_ ( .A(\EXU/_0232_ ), .Z(\EXU/_1526_ ) );
BUF_X1 \EXU/_3182_ ( .A(\_IDU_io_out_bits_rd1 [31] ), .Z(\EXU/_0703_ ) );
BUF_X1 \EXU/_3183_ ( .A(\EXU/_0233_ ), .Z(\EXU/_1527_ ) );
BUF_X1 \EXU/_3184_ ( .A(\_IDU_io_out_bits_rd2 [0] ), .Z(\EXU/_0711_ ) );
BUF_X1 \EXU/_3185_ ( .A(\EXU/_0234_ ), .Z(\EXU/_1528_ ) );
BUF_X1 \EXU/_3186_ ( .A(\_IDU_io_out_bits_rd2 [1] ), .Z(\EXU/_0722_ ) );
BUF_X1 \EXU/_3187_ ( .A(\EXU/_0235_ ), .Z(\EXU/_1529_ ) );
BUF_X1 \EXU/_3188_ ( .A(\_IDU_io_out_bits_rd2 [2] ), .Z(\EXU/_0733_ ) );
BUF_X1 \EXU/_3189_ ( .A(\EXU/_0236_ ), .Z(\EXU/_1530_ ) );
BUF_X1 \EXU/_3190_ ( .A(\_IDU_io_out_bits_rd2 [3] ), .Z(\EXU/_0736_ ) );
BUF_X1 \EXU/_3191_ ( .A(\EXU/_0237_ ), .Z(\EXU/_1531_ ) );
BUF_X1 \EXU/_3192_ ( .A(\_IDU_io_out_bits_rd2 [4] ), .Z(\EXU/_0737_ ) );
BUF_X1 \EXU/_3193_ ( .A(\EXU/_0238_ ), .Z(\EXU/_1532_ ) );
BUF_X1 \EXU/_3194_ ( .A(\_IDU_io_out_bits_rd2 [5] ), .Z(\EXU/_0738_ ) );
BUF_X1 \EXU/_3195_ ( .A(\EXU/_0239_ ), .Z(\EXU/_1533_ ) );
BUF_X1 \EXU/_3196_ ( .A(\_IDU_io_out_bits_rd2 [6] ), .Z(\EXU/_0739_ ) );
BUF_X1 \EXU/_3197_ ( .A(\EXU/_0240_ ), .Z(\EXU/_1534_ ) );
BUF_X1 \EXU/_3198_ ( .A(\_IDU_io_out_bits_rd2 [7] ), .Z(\EXU/_0740_ ) );
BUF_X1 \EXU/_3199_ ( .A(\EXU/_0241_ ), .Z(\EXU/_1535_ ) );
BUF_X1 \EXU/_3200_ ( .A(\_IDU_io_out_bits_rd2 [8] ), .Z(\EXU/_0741_ ) );
BUF_X1 \EXU/_3201_ ( .A(\EXU/_0242_ ), .Z(\EXU/_1536_ ) );
BUF_X1 \EXU/_3202_ ( .A(\_IDU_io_out_bits_rd2 [9] ), .Z(\EXU/_0742_ ) );
BUF_X1 \EXU/_3203_ ( .A(\EXU/_0243_ ), .Z(\EXU/_1537_ ) );
BUF_X1 \EXU/_3204_ ( .A(\_IDU_io_out_bits_rd2 [10] ), .Z(\EXU/_0712_ ) );
BUF_X1 \EXU/_3205_ ( .A(\EXU/_0244_ ), .Z(\EXU/_1538_ ) );
BUF_X1 \EXU/_3206_ ( .A(\_IDU_io_out_bits_rd2 [11] ), .Z(\EXU/_0713_ ) );
BUF_X1 \EXU/_3207_ ( .A(\EXU/_0245_ ), .Z(\EXU/_1539_ ) );
BUF_X1 \EXU/_3208_ ( .A(\_IDU_io_out_bits_rd2 [12] ), .Z(\EXU/_0714_ ) );
BUF_X1 \EXU/_3209_ ( .A(\EXU/_0246_ ), .Z(\EXU/_1540_ ) );
BUF_X1 \EXU/_3210_ ( .A(\_IDU_io_out_bits_rd2 [13] ), .Z(\EXU/_0715_ ) );
BUF_X1 \EXU/_3211_ ( .A(\EXU/_0247_ ), .Z(\EXU/_1541_ ) );
BUF_X1 \EXU/_3212_ ( .A(\_IDU_io_out_bits_rd2 [14] ), .Z(\EXU/_0716_ ) );
BUF_X1 \EXU/_3213_ ( .A(\EXU/_0248_ ), .Z(\EXU/_1542_ ) );
BUF_X1 \EXU/_3214_ ( .A(\_IDU_io_out_bits_rd2 [15] ), .Z(\EXU/_0717_ ) );
BUF_X1 \EXU/_3215_ ( .A(\EXU/_0249_ ), .Z(\EXU/_1543_ ) );
BUF_X1 \EXU/_3216_ ( .A(\_IDU_io_out_bits_rd2 [16] ), .Z(\EXU/_0718_ ) );
BUF_X1 \EXU/_3217_ ( .A(\EXU/_0250_ ), .Z(\EXU/_1544_ ) );
BUF_X1 \EXU/_3218_ ( .A(\_IDU_io_out_bits_rd2 [17] ), .Z(\EXU/_0719_ ) );
BUF_X1 \EXU/_3219_ ( .A(\EXU/_0251_ ), .Z(\EXU/_1545_ ) );
BUF_X1 \EXU/_3220_ ( .A(\_IDU_io_out_bits_rd2 [18] ), .Z(\EXU/_0720_ ) );
BUF_X1 \EXU/_3221_ ( .A(\EXU/_0252_ ), .Z(\EXU/_1546_ ) );
BUF_X1 \EXU/_3222_ ( .A(\_IDU_io_out_bits_rd2 [19] ), .Z(\EXU/_0721_ ) );
BUF_X1 \EXU/_3223_ ( .A(\EXU/_0253_ ), .Z(\EXU/_1547_ ) );
BUF_X1 \EXU/_3224_ ( .A(\_IDU_io_out_bits_rd2 [20] ), .Z(\EXU/_0723_ ) );
BUF_X1 \EXU/_3225_ ( .A(\EXU/_0254_ ), .Z(\EXU/_1548_ ) );
BUF_X1 \EXU/_3226_ ( .A(\_IDU_io_out_bits_rd2 [21] ), .Z(\EXU/_0724_ ) );
BUF_X1 \EXU/_3227_ ( .A(\EXU/_0255_ ), .Z(\EXU/_1549_ ) );
BUF_X1 \EXU/_3228_ ( .A(\_IDU_io_out_bits_rd2 [22] ), .Z(\EXU/_0725_ ) );
BUF_X1 \EXU/_3229_ ( .A(\EXU/_0256_ ), .Z(\EXU/_1550_ ) );
BUF_X1 \EXU/_3230_ ( .A(\_IDU_io_out_bits_rd2 [23] ), .Z(\EXU/_0726_ ) );
BUF_X1 \EXU/_3231_ ( .A(\EXU/_0257_ ), .Z(\EXU/_1551_ ) );
BUF_X1 \EXU/_3232_ ( .A(\_IDU_io_out_bits_rd2 [24] ), .Z(\EXU/_0727_ ) );
BUF_X1 \EXU/_3233_ ( .A(\EXU/_0258_ ), .Z(\EXU/_1552_ ) );
BUF_X1 \EXU/_3234_ ( .A(\_IDU_io_out_bits_rd2 [25] ), .Z(\EXU/_0728_ ) );
BUF_X1 \EXU/_3235_ ( .A(\EXU/_0259_ ), .Z(\EXU/_1553_ ) );
BUF_X1 \EXU/_3236_ ( .A(\_IDU_io_out_bits_rd2 [26] ), .Z(\EXU/_0729_ ) );
BUF_X1 \EXU/_3237_ ( .A(\EXU/_0260_ ), .Z(\EXU/_1554_ ) );
BUF_X1 \EXU/_3238_ ( .A(\_IDU_io_out_bits_rd2 [27] ), .Z(\EXU/_0730_ ) );
BUF_X1 \EXU/_3239_ ( .A(\EXU/_0261_ ), .Z(\EXU/_1555_ ) );
BUF_X1 \EXU/_3240_ ( .A(\_IDU_io_out_bits_rd2 [28] ), .Z(\EXU/_0731_ ) );
BUF_X1 \EXU/_3241_ ( .A(\EXU/_0262_ ), .Z(\EXU/_1556_ ) );
BUF_X1 \EXU/_3242_ ( .A(\_IDU_io_out_bits_rd2 [29] ), .Z(\EXU/_0732_ ) );
BUF_X1 \EXU/_3243_ ( .A(\EXU/_0263_ ), .Z(\EXU/_1557_ ) );
BUF_X1 \EXU/_3244_ ( .A(\_IDU_io_out_bits_rd2 [30] ), .Z(\EXU/_0734_ ) );
BUF_X1 \EXU/_3245_ ( .A(\EXU/_0264_ ), .Z(\EXU/_1558_ ) );
BUF_X1 \EXU/_3246_ ( .A(\_IDU_io_out_bits_rd2 [31] ), .Z(\EXU/_0735_ ) );
BUF_X1 \EXU/_3247_ ( .A(\EXU/_0265_ ), .Z(\EXU/_1559_ ) );
BUF_X1 \EXU/_3248_ ( .A(\_IDU_io_out_bits_imm [0] ), .Z(\EXU/_0615_ ) );
BUF_X1 \EXU/_3249_ ( .A(\EXU/_0266_ ), .Z(\EXU/_1560_ ) );
BUF_X1 \EXU/_3250_ ( .A(\_IDU_io_out_bits_imm [1] ), .Z(\EXU/_0626_ ) );
BUF_X1 \EXU/_3251_ ( .A(\EXU/_0267_ ), .Z(\EXU/_1561_ ) );
BUF_X1 \EXU/_3252_ ( .A(\_IDU_io_out_bits_imm [2] ), .Z(\EXU/_0637_ ) );
BUF_X1 \EXU/_3253_ ( .A(\EXU/_0268_ ), .Z(\EXU/_1562_ ) );
BUF_X1 \EXU/_3254_ ( .A(\_IDU_io_out_bits_imm [3] ), .Z(\EXU/_0640_ ) );
BUF_X1 \EXU/_3255_ ( .A(\EXU/_0269_ ), .Z(\EXU/_1563_ ) );
BUF_X1 \EXU/_3256_ ( .A(\_IDU_io_out_bits_imm [4] ), .Z(\EXU/_0641_ ) );
BUF_X1 \EXU/_3257_ ( .A(\EXU/_0270_ ), .Z(\EXU/_1564_ ) );
BUF_X1 \EXU/_3258_ ( .A(\_IDU_io_out_bits_imm [5] ), .Z(\EXU/_0642_ ) );
BUF_X1 \EXU/_3259_ ( .A(\EXU/_0271_ ), .Z(\EXU/_1565_ ) );
BUF_X1 \EXU/_3260_ ( .A(\_IDU_io_out_bits_imm [6] ), .Z(\EXU/_0643_ ) );
BUF_X1 \EXU/_3261_ ( .A(\EXU/_0272_ ), .Z(\EXU/_1566_ ) );
BUF_X1 \EXU/_3262_ ( .A(\_IDU_io_out_bits_imm [7] ), .Z(\EXU/_0644_ ) );
BUF_X1 \EXU/_3263_ ( .A(\EXU/_0273_ ), .Z(\EXU/_1567_ ) );
BUF_X1 \EXU/_3264_ ( .A(\_IDU_io_out_bits_imm [8] ), .Z(\EXU/_0645_ ) );
BUF_X1 \EXU/_3265_ ( .A(\EXU/_0274_ ), .Z(\EXU/_1568_ ) );
BUF_X1 \EXU/_3266_ ( .A(\_IDU_io_out_bits_imm [9] ), .Z(\EXU/_0646_ ) );
BUF_X1 \EXU/_3267_ ( .A(\EXU/_0275_ ), .Z(\EXU/_1569_ ) );
BUF_X1 \EXU/_3268_ ( .A(\_IDU_io_out_bits_imm [10] ), .Z(\EXU/_0616_ ) );
BUF_X1 \EXU/_3269_ ( .A(\EXU/_0276_ ), .Z(\EXU/_1570_ ) );
BUF_X1 \EXU/_3270_ ( .A(\_IDU_io_out_bits_imm [11] ), .Z(\EXU/_0617_ ) );
BUF_X1 \EXU/_3271_ ( .A(\EXU/_0277_ ), .Z(\EXU/_1571_ ) );
BUF_X1 \EXU/_3272_ ( .A(\_IDU_io_out_bits_imm [12] ), .Z(\EXU/_0618_ ) );
BUF_X1 \EXU/_3273_ ( .A(\EXU/_0278_ ), .Z(\EXU/_1572_ ) );
BUF_X1 \EXU/_3274_ ( .A(\_IDU_io_out_bits_imm [13] ), .Z(\EXU/_0619_ ) );
BUF_X1 \EXU/_3275_ ( .A(\EXU/_0279_ ), .Z(\EXU/_1573_ ) );
BUF_X1 \EXU/_3276_ ( .A(\_IDU_io_out_bits_imm [14] ), .Z(\EXU/_0620_ ) );
BUF_X1 \EXU/_3277_ ( .A(\EXU/_0280_ ), .Z(\EXU/_1574_ ) );
BUF_X1 \EXU/_3278_ ( .A(\_IDU_io_out_bits_imm [15] ), .Z(\EXU/_0621_ ) );
BUF_X1 \EXU/_3279_ ( .A(\EXU/_0281_ ), .Z(\EXU/_1575_ ) );
BUF_X1 \EXU/_3280_ ( .A(\_IDU_io_out_bits_imm [16] ), .Z(\EXU/_0622_ ) );
BUF_X1 \EXU/_3281_ ( .A(\EXU/_0282_ ), .Z(\EXU/_1576_ ) );
BUF_X1 \EXU/_3282_ ( .A(\_IDU_io_out_bits_imm [17] ), .Z(\EXU/_0623_ ) );
BUF_X1 \EXU/_3283_ ( .A(\EXU/_0283_ ), .Z(\EXU/_1577_ ) );
BUF_X1 \EXU/_3284_ ( .A(\_IDU_io_out_bits_imm [18] ), .Z(\EXU/_0624_ ) );
BUF_X1 \EXU/_3285_ ( .A(\EXU/_0284_ ), .Z(\EXU/_1578_ ) );
BUF_X1 \EXU/_3286_ ( .A(\_IDU_io_out_bits_imm [19] ), .Z(\EXU/_0625_ ) );
BUF_X1 \EXU/_3287_ ( .A(\EXU/_0285_ ), .Z(\EXU/_1579_ ) );
BUF_X1 \EXU/_3288_ ( .A(\_IDU_io_out_bits_imm [20] ), .Z(\EXU/_0627_ ) );
BUF_X1 \EXU/_3289_ ( .A(\EXU/_0286_ ), .Z(\EXU/_1580_ ) );
BUF_X1 \EXU/_3290_ ( .A(\_IDU_io_out_bits_imm [21] ), .Z(\EXU/_0628_ ) );
BUF_X1 \EXU/_3291_ ( .A(\EXU/_0287_ ), .Z(\EXU/_1581_ ) );
BUF_X1 \EXU/_3292_ ( .A(\_IDU_io_out_bits_imm [22] ), .Z(\EXU/_0629_ ) );
BUF_X1 \EXU/_3293_ ( .A(\EXU/_0288_ ), .Z(\EXU/_1582_ ) );
BUF_X1 \EXU/_3294_ ( .A(\_IDU_io_out_bits_imm [23] ), .Z(\EXU/_0630_ ) );
BUF_X1 \EXU/_3295_ ( .A(\EXU/_0289_ ), .Z(\EXU/_1583_ ) );
BUF_X1 \EXU/_3296_ ( .A(\_IDU_io_out_bits_imm [24] ), .Z(\EXU/_0631_ ) );
BUF_X1 \EXU/_3297_ ( .A(\EXU/_0290_ ), .Z(\EXU/_1584_ ) );
BUF_X1 \EXU/_3298_ ( .A(\_IDU_io_out_bits_imm [25] ), .Z(\EXU/_0632_ ) );
BUF_X1 \EXU/_3299_ ( .A(\EXU/_0291_ ), .Z(\EXU/_1585_ ) );
BUF_X1 \EXU/_3300_ ( .A(\_IDU_io_out_bits_imm [26] ), .Z(\EXU/_0633_ ) );
BUF_X1 \EXU/_3301_ ( .A(\EXU/_0292_ ), .Z(\EXU/_1586_ ) );
BUF_X1 \EXU/_3302_ ( .A(\_IDU_io_out_bits_imm [27] ), .Z(\EXU/_0634_ ) );
BUF_X1 \EXU/_3303_ ( .A(\EXU/_0293_ ), .Z(\EXU/_1587_ ) );
BUF_X1 \EXU/_3304_ ( .A(\_IDU_io_out_bits_imm [28] ), .Z(\EXU/_0635_ ) );
BUF_X1 \EXU/_3305_ ( .A(\EXU/_0294_ ), .Z(\EXU/_1588_ ) );
BUF_X1 \EXU/_3306_ ( .A(\_IDU_io_out_bits_imm [29] ), .Z(\EXU/_0636_ ) );
BUF_X1 \EXU/_3307_ ( .A(\EXU/_0295_ ), .Z(\EXU/_1589_ ) );
BUF_X1 \EXU/_3308_ ( .A(\_IDU_io_out_bits_imm [30] ), .Z(\EXU/_0638_ ) );
BUF_X1 \EXU/_3309_ ( .A(\EXU/_0296_ ), .Z(\EXU/_1590_ ) );
BUF_X1 \EXU/_3310_ ( .A(\_IDU_io_out_bits_imm [31] ), .Z(\EXU/_0639_ ) );
BUF_X1 \EXU/_3311_ ( .A(\EXU/_0297_ ), .Z(\EXU/_1591_ ) );
BUF_X1 \EXU/_3312_ ( .A(\_IDU_io_out_bits_uimm [0] ), .Z(\EXU/_0743_ ) );
BUF_X1 \EXU/_3313_ ( .A(\EXU/_0298_ ), .Z(\EXU/_1592_ ) );
BUF_X1 \EXU/_3314_ ( .A(\_IDU_io_out_bits_uimm [1] ), .Z(\EXU/_0754_ ) );
BUF_X1 \EXU/_3315_ ( .A(\EXU/_0299_ ), .Z(\EXU/_1593_ ) );
BUF_X1 \EXU/_3316_ ( .A(\_IDU_io_out_bits_uimm [2] ), .Z(\EXU/_0765_ ) );
BUF_X1 \EXU/_3317_ ( .A(\EXU/_0300_ ), .Z(\EXU/_1594_ ) );
BUF_X1 \EXU/_3318_ ( .A(\_IDU_io_out_bits_uimm [3] ), .Z(\EXU/_0768_ ) );
BUF_X1 \EXU/_3319_ ( .A(\EXU/_0301_ ), .Z(\EXU/_1595_ ) );
BUF_X1 \EXU/_3320_ ( .A(\_IDU_io_out_bits_uimm [4] ), .Z(\EXU/_0769_ ) );
BUF_X1 \EXU/_3321_ ( .A(\EXU/_0302_ ), .Z(\EXU/_1596_ ) );
BUF_X1 \EXU/_3322_ ( .A(\_IDU_io_out_bits_uimm [5] ), .Z(\EXU/_0770_ ) );
BUF_X1 \EXU/_3323_ ( .A(\EXU/_0303_ ), .Z(\EXU/_1597_ ) );
BUF_X1 \EXU/_3324_ ( .A(\_IDU_io_out_bits_uimm [6] ), .Z(\EXU/_0771_ ) );
BUF_X1 \EXU/_3325_ ( .A(\EXU/_0304_ ), .Z(\EXU/_1598_ ) );
BUF_X1 \EXU/_3326_ ( .A(\_IDU_io_out_bits_uimm [7] ), .Z(\EXU/_0772_ ) );
BUF_X1 \EXU/_3327_ ( .A(\EXU/_0305_ ), .Z(\EXU/_1599_ ) );
BUF_X1 \EXU/_3328_ ( .A(\_IDU_io_out_bits_uimm [8] ), .Z(\EXU/_0773_ ) );
BUF_X1 \EXU/_3329_ ( .A(\EXU/_0306_ ), .Z(\EXU/_1600_ ) );
BUF_X1 \EXU/_3330_ ( .A(\_IDU_io_out_bits_uimm [9] ), .Z(\EXU/_0774_ ) );
BUF_X1 \EXU/_3331_ ( .A(\EXU/_0307_ ), .Z(\EXU/_1601_ ) );
BUF_X1 \EXU/_3332_ ( .A(\_IDU_io_out_bits_uimm [10] ), .Z(\EXU/_0744_ ) );
BUF_X1 \EXU/_3333_ ( .A(\EXU/_0308_ ), .Z(\EXU/_1602_ ) );
BUF_X1 \EXU/_3334_ ( .A(\_IDU_io_out_bits_uimm [11] ), .Z(\EXU/_0745_ ) );
BUF_X1 \EXU/_3335_ ( .A(\EXU/_0309_ ), .Z(\EXU/_1603_ ) );
BUF_X1 \EXU/_3336_ ( .A(\_IDU_io_out_bits_uimm [12] ), .Z(\EXU/_0746_ ) );
BUF_X1 \EXU/_3337_ ( .A(\EXU/_0310_ ), .Z(\EXU/_1604_ ) );
BUF_X1 \EXU/_3338_ ( .A(\_IDU_io_out_bits_uimm [13] ), .Z(\EXU/_0747_ ) );
BUF_X1 \EXU/_3339_ ( .A(\EXU/_0311_ ), .Z(\EXU/_1605_ ) );
BUF_X1 \EXU/_3340_ ( .A(\_IDU_io_out_bits_uimm [14] ), .Z(\EXU/_0748_ ) );
BUF_X1 \EXU/_3341_ ( .A(\EXU/_0312_ ), .Z(\EXU/_1606_ ) );
BUF_X1 \EXU/_3342_ ( .A(\_IDU_io_out_bits_uimm [15] ), .Z(\EXU/_0749_ ) );
BUF_X1 \EXU/_3343_ ( .A(\EXU/_0313_ ), .Z(\EXU/_1607_ ) );
BUF_X1 \EXU/_3344_ ( .A(\_IDU_io_out_bits_uimm [16] ), .Z(\EXU/_0750_ ) );
BUF_X1 \EXU/_3345_ ( .A(\EXU/_0314_ ), .Z(\EXU/_1608_ ) );
BUF_X1 \EXU/_3346_ ( .A(\_IDU_io_out_bits_uimm [17] ), .Z(\EXU/_0751_ ) );
BUF_X1 \EXU/_3347_ ( .A(\EXU/_0315_ ), .Z(\EXU/_1609_ ) );
BUF_X1 \EXU/_3348_ ( .A(\_IDU_io_out_bits_uimm [18] ), .Z(\EXU/_0752_ ) );
BUF_X1 \EXU/_3349_ ( .A(\EXU/_0316_ ), .Z(\EXU/_1610_ ) );
BUF_X1 \EXU/_3350_ ( .A(\_IDU_io_out_bits_uimm [19] ), .Z(\EXU/_0753_ ) );
BUF_X1 \EXU/_3351_ ( .A(\EXU/_0317_ ), .Z(\EXU/_1611_ ) );
BUF_X1 \EXU/_3352_ ( .A(\_IDU_io_out_bits_uimm [20] ), .Z(\EXU/_0755_ ) );
BUF_X1 \EXU/_3353_ ( .A(\EXU/_0318_ ), .Z(\EXU/_1612_ ) );
BUF_X1 \EXU/_3354_ ( .A(\_IDU_io_out_bits_uimm [21] ), .Z(\EXU/_0756_ ) );
BUF_X1 \EXU/_3355_ ( .A(\EXU/_0319_ ), .Z(\EXU/_1613_ ) );
BUF_X1 \EXU/_3356_ ( .A(\_IDU_io_out_bits_uimm [22] ), .Z(\EXU/_0757_ ) );
BUF_X1 \EXU/_3357_ ( .A(\EXU/_0320_ ), .Z(\EXU/_1614_ ) );
BUF_X1 \EXU/_3358_ ( .A(\_IDU_io_out_bits_uimm [23] ), .Z(\EXU/_0758_ ) );
BUF_X1 \EXU/_3359_ ( .A(\EXU/_0321_ ), .Z(\EXU/_1615_ ) );
BUF_X1 \EXU/_3360_ ( .A(\_IDU_io_out_bits_uimm [24] ), .Z(\EXU/_0759_ ) );
BUF_X1 \EXU/_3361_ ( .A(\EXU/_0322_ ), .Z(\EXU/_1616_ ) );
BUF_X1 \EXU/_3362_ ( .A(\_IDU_io_out_bits_uimm [25] ), .Z(\EXU/_0760_ ) );
BUF_X1 \EXU/_3363_ ( .A(\EXU/_0323_ ), .Z(\EXU/_1617_ ) );
BUF_X1 \EXU/_3364_ ( .A(\_IDU_io_out_bits_uimm [26] ), .Z(\EXU/_0761_ ) );
BUF_X1 \EXU/_3365_ ( .A(\EXU/_0324_ ), .Z(\EXU/_1618_ ) );
BUF_X1 \EXU/_3366_ ( .A(\_IDU_io_out_bits_uimm [27] ), .Z(\EXU/_0762_ ) );
BUF_X1 \EXU/_3367_ ( .A(\EXU/_0325_ ), .Z(\EXU/_1619_ ) );
BUF_X1 \EXU/_3368_ ( .A(\_IDU_io_out_bits_uimm [28] ), .Z(\EXU/_0763_ ) );
BUF_X1 \EXU/_3369_ ( .A(\EXU/_0326_ ), .Z(\EXU/_1620_ ) );
BUF_X1 \EXU/_3370_ ( .A(\_IDU_io_out_bits_uimm [29] ), .Z(\EXU/_0764_ ) );
BUF_X1 \EXU/_3371_ ( .A(\EXU/_0327_ ), .Z(\EXU/_1621_ ) );
BUF_X1 \EXU/_3372_ ( .A(\_IDU_io_out_bits_uimm [30] ), .Z(\EXU/_0766_ ) );
BUF_X1 \EXU/_3373_ ( .A(\EXU/_0328_ ), .Z(\EXU/_1622_ ) );
BUF_X1 \EXU/_3374_ ( .A(\_IDU_io_out_bits_uimm [31] ), .Z(\EXU/_0767_ ) );
BUF_X1 \EXU/_3375_ ( .A(\EXU/_0329_ ), .Z(\EXU/_1623_ ) );
BUF_X1 \EXU/_3376_ ( .A(_IDU_io_out_bits_control_aluASrc ), .Z(\EXU/_0596_ ) );
BUF_X1 \EXU/_3377_ ( .A(\EXU/_0330_ ), .Z(\EXU/_1624_ ) );
BUF_X1 \EXU/_3378_ ( .A(\_IDU_io_out_bits_control_aluBSrc [0] ), .Z(\EXU/_0597_ ) );
BUF_X1 \EXU/_3379_ ( .A(\EXU/_0331_ ), .Z(\EXU/_1625_ ) );
BUF_X1 \EXU/_3380_ ( .A(\_IDU_io_out_bits_control_aluBSrc [1] ), .Z(\EXU/_0598_ ) );
BUF_X1 \EXU/_3381_ ( .A(\EXU/_0332_ ), .Z(\EXU/_1626_ ) );
BUF_X1 \EXU/_3382_ ( .A(\EXU/in_control_aluCtr [0] ), .Z(\EXU/_0384_ ) );
BUF_X1 \EXU/_3383_ ( .A(\_IDU_io_out_bits_control_aluCtr [0] ), .Z(\EXU/_0599_ ) );
BUF_X1 \EXU/_3384_ ( .A(\EXU/_0333_ ), .Z(\EXU/_1627_ ) );
BUF_X1 \EXU/_3385_ ( .A(\EXU/in_control_aluCtr [1] ), .Z(\EXU/_0385_ ) );
BUF_X1 \EXU/_3386_ ( .A(\_IDU_io_out_bits_control_aluCtr [1] ), .Z(\EXU/_0600_ ) );
BUF_X1 \EXU/_3387_ ( .A(\EXU/_0334_ ), .Z(\EXU/_1628_ ) );
BUF_X1 \EXU/_3388_ ( .A(\EXU/in_control_aluCtr [2] ), .Z(\EXU/_0386_ ) );
BUF_X1 \EXU/_3389_ ( .A(\_IDU_io_out_bits_control_aluCtr [2] ), .Z(\EXU/_0601_ ) );
BUF_X1 \EXU/_3390_ ( .A(\EXU/_0335_ ), .Z(\EXU/_1629_ ) );
BUF_X1 \EXU/_3391_ ( .A(\EXU/in_control_aluCtr [3] ), .Z(\EXU/_0387_ ) );
BUF_X1 \EXU/_3392_ ( .A(\_IDU_io_out_bits_control_aluCtr [3] ), .Z(\EXU/_0602_ ) );
BUF_X1 \EXU/_3393_ ( .A(\EXU/_0336_ ), .Z(\EXU/_1630_ ) );
BUF_X1 \EXU/_3394_ ( .A(_IDU_io_out_bits_control_csrSrc ), .Z(\EXU/_0609_ ) );
BUF_X1 \EXU/_3395_ ( .A(\EXU/_0337_ ), .Z(\EXU/_1631_ ) );
BUF_X1 \EXU/_3396_ ( .A(\_IDU_io_out_bits_control_csrCtr [0] ), .Z(\EXU/_0606_ ) );
BUF_X1 \EXU/_3397_ ( .A(\EXU/_0338_ ), .Z(\EXU/_1632_ ) );
BUF_X1 \EXU/_3398_ ( .A(\_IDU_io_out_bits_control_csrCtr [1] ), .Z(\EXU/_0607_ ) );
BUF_X1 \EXU/_3399_ ( .A(\EXU/_0339_ ), .Z(\EXU/_1633_ ) );
BUF_X1 \EXU/_3400_ ( .A(\_IDU_io_out_bits_control_csrCtr [2] ), .Z(\EXU/_0608_ ) );
BUF_X1 \EXU/_3401_ ( .A(\EXU/_0340_ ), .Z(\EXU/_1634_ ) );
BUF_X1 \EXU/_3402_ ( .A(\EXU/in_control_brType [0] ), .Z(\EXU/_0388_ ) );
BUF_X1 \EXU/_3403_ ( .A(\_IDU_io_out_bits_control_brType [0] ), .Z(\EXU/_0603_ ) );
BUF_X1 \EXU/_3404_ ( .A(\EXU/_0341_ ), .Z(\EXU/_1635_ ) );
BUF_X1 \EXU/_3405_ ( .A(\EXU/in_control_brType [1] ), .Z(\EXU/_0389_ ) );
BUF_X1 \EXU/_3406_ ( .A(\_IDU_io_out_bits_control_brType [1] ), .Z(\EXU/_0604_ ) );
BUF_X1 \EXU/_3407_ ( .A(\EXU/_0342_ ), .Z(\EXU/_1636_ ) );
BUF_X1 \EXU/_3408_ ( .A(\EXU/in_control_brType [2] ), .Z(\EXU/_0390_ ) );
BUF_X1 \EXU/_3409_ ( .A(\_IDU_io_out_bits_control_brType [2] ), .Z(\EXU/_0605_ ) );
BUF_X1 \EXU/_3410_ ( .A(\EXU/_0343_ ), .Z(\EXU/_1637_ ) );
BUF_X1 \EXU/_3411_ ( .A(_EXU_io_LSUIn_bits_ren ), .Z(\EXU/_0526_ ) );
BUF_X1 \EXU/_3412_ ( .A(\EXU/_0344_ ), .Z(\EXU/_1638_ ) );
BUF_X1 \EXU/_3413_ ( .A(_EXU_io_LSUIn_bits_wen ), .Z(\EXU/_0559_ ) );
BUF_X1 \EXU/_3414_ ( .A(\EXU/_0345_ ), .Z(\EXU/_1639_ ) );
BUF_X1 \EXU/_3415_ ( .A(\_EXU_io_LSUIn_bits_memOp [0] ), .Z(\EXU/_0523_ ) );
BUF_X1 \EXU/_3416_ ( .A(\_IDU_io_out_bits_control_memOp [0] ), .Z(\EXU/_0610_ ) );
BUF_X1 \EXU/_3417_ ( .A(\EXU/_0346_ ), .Z(\EXU/_1640_ ) );
BUF_X1 \EXU/_3418_ ( .A(\_EXU_io_LSUIn_bits_memOp [1] ), .Z(\EXU/_0524_ ) );
BUF_X1 \EXU/_3419_ ( .A(\_IDU_io_out_bits_control_memOp [1] ), .Z(\EXU/_0611_ ) );
BUF_X1 \EXU/_3420_ ( .A(\EXU/_0347_ ), .Z(\EXU/_1641_ ) );
BUF_X1 \EXU/_3421_ ( .A(\_EXU_io_LSUIn_bits_memOp [2] ), .Z(\EXU/_0525_ ) );
BUF_X1 \EXU/_3422_ ( .A(\_IDU_io_out_bits_control_memOp [2] ), .Z(\EXU/_0612_ ) );
BUF_X1 \EXU/_3423_ ( .A(\EXU/_0348_ ), .Z(\EXU/_1642_ ) );
BUF_X1 \EXU/_3424_ ( .A(reset ), .Z(\EXU/_1214_ ) );
BUF_X1 \EXU/_3425_ ( .A(\EXU/_0168_ ), .Z(\EXU/_1462_ ) );
BUF_X1 \EXU/_3426_ ( .A(\EXU/_0169_ ), .Z(\EXU/_1463_ ) );
XOR2_X1 \EXU/ALU/_458_ ( .A(\EXU/ALU/_026_ ), .B(\EXU/ALU/_001_ ), .Z(\EXU/ALU/_168_ ) );
OR2_X1 \EXU/ALU/_459_ ( .A1(\EXU/ALU/_168_ ), .A2(\EXU/ALU/_038_ ), .ZN(\EXU/ALU/_169_ ) );
XNOR2_X1 \EXU/ALU/_460_ ( .A(\EXU/ALU/_037_ ), .B(\EXU/ALU/_000_ ), .ZN(\EXU/ALU/_170_ ) );
NAND2_X1 \EXU/ALU/_461_ ( .A1(\EXU/ALU/_170_ ), .A2(\EXU/ALU/_038_ ), .ZN(\EXU/ALU/_171_ ) );
AND2_X1 \EXU/ALU/_462_ ( .A1(\EXU/ALU/_169_ ), .A2(\EXU/ALU/_171_ ), .ZN(\EXU/ALU/_167_ ) );
INV_X4 \EXU/ALU/_463_ ( .A(fanout_net_12 ), .ZN(\EXU/ALU/_172_ ) );
INV_X32 \EXU/ALU/_464_ ( .A(fanout_net_14 ), .ZN(\EXU/ALU/_173_ ) );
BUF_X4 \EXU/ALU/_465_ ( .A(\EXU/ALU/_173_ ), .Z(\EXU/ALU/_174_ ) );
AND3_X1 \EXU/ALU/_466_ ( .A1(\EXU/ALU/_172_ ), .A2(\EXU/ALU/_174_ ), .A3(fanout_net_13 ), .ZN(\EXU/ALU/_175_ ) );
NAND3_X1 \EXU/ALU/_467_ ( .A1(\EXU/ALU/_169_ ), .A2(\EXU/ALU/_171_ ), .A3(\EXU/ALU/_175_ ), .ZN(\EXU/ALU/_176_ ) );
OR2_X1 \EXU/ALU/_468_ ( .A1(\EXU/ALU/_135_ ), .A2(\EXU/ALU/_103_ ), .ZN(\EXU/ALU/_177_ ) );
NOR2_X4 \EXU/ALU/_469_ ( .A1(fanout_net_12 ), .A2(fanout_net_13 ), .ZN(\EXU/ALU/_178_ ) );
NAND2_X1 \EXU/ALU/_470_ ( .A1(\EXU/ALU/_135_ ), .A2(\EXU/ALU/_103_ ), .ZN(\EXU/ALU/_179_ ) );
AND3_X1 \EXU/ALU/_471_ ( .A1(\EXU/ALU/_178_ ), .A2(fanout_net_14 ), .A3(\EXU/ALU/_179_ ), .ZN(\EXU/ALU/_180_ ) );
NAND2_X1 \EXU/ALU/_472_ ( .A1(\EXU/ALU/_172_ ), .A2(fanout_net_13 ), .ZN(\EXU/ALU/_181_ ) );
NOR2_X2 \EXU/ALU/_473_ ( .A1(\EXU/ALU/_181_ ), .A2(\EXU/ALU/_173_ ), .ZN(\EXU/ALU/_182_ ) );
BUF_X4 \EXU/ALU/_474_ ( .A(\EXU/ALU/_182_ ), .Z(\EXU/ALU/_183_ ) );
OAI21_X1 \EXU/ALU/_475_ ( .A(\EXU/ALU/_177_ ), .B1(\EXU/ALU/_180_ ), .B2(\EXU/ALU/_183_ ), .ZN(\EXU/ALU/_184_ ) );
AND2_X2 \EXU/ALU/_476_ ( .A1(fanout_net_12 ), .A2(fanout_net_13 ), .ZN(\EXU/ALU/_185_ ) );
BUF_X4 \EXU/ALU/_477_ ( .A(\EXU/ALU/_173_ ), .Z(\EXU/ALU/_186_ ) );
OAI211_X2 \EXU/ALU/_478_ ( .A(\EXU/ALU/_185_ ), .B(\EXU/ALU/_135_ ), .C1(\EXU/ALU/_103_ ), .C2(\EXU/ALU/_186_ ), .ZN(\EXU/ALU/_187_ ) );
AND3_X1 \EXU/ALU/_479_ ( .A1(\EXU/ALU/_178_ ), .A2(\EXU/ALU/_174_ ), .A3(\EXU/ALU/_002_ ), .ZN(\EXU/ALU/_188_ ) );
NOR2_X2 \EXU/ALU/_480_ ( .A1(\EXU/ALU/_172_ ), .A2(fanout_net_13 ), .ZN(\EXU/ALU/_189_ ) );
BUF_X4 \EXU/ALU/_481_ ( .A(\EXU/ALU/_189_ ), .Z(\EXU/ALU/_190_ ) );
AOI21_X1 \EXU/ALU/_482_ ( .A(\EXU/ALU/_188_ ), .B1(\EXU/ALU/_039_ ), .B2(\EXU/ALU/_190_ ), .ZN(\EXU/ALU/_191_ ) );
NAND4_X1 \EXU/ALU/_483_ ( .A1(\EXU/ALU/_176_ ), .A2(\EXU/ALU/_184_ ), .A3(\EXU/ALU/_187_ ), .A4(\EXU/ALU/_191_ ), .ZN(\EXU/ALU/_071_ ) );
OR2_X1 \EXU/ALU/_484_ ( .A1(\EXU/ALU/_146_ ), .A2(\EXU/ALU/_114_ ), .ZN(\EXU/ALU/_192_ ) );
BUF_X4 \EXU/ALU/_485_ ( .A(\EXU/ALU/_178_ ), .Z(\EXU/ALU/_193_ ) );
NAND2_X1 \EXU/ALU/_486_ ( .A1(\EXU/ALU/_146_ ), .A2(\EXU/ALU/_114_ ), .ZN(\EXU/ALU/_194_ ) );
NAND4_X1 \EXU/ALU/_487_ ( .A1(\EXU/ALU/_192_ ), .A2(fanout_net_14 ), .A3(\EXU/ALU/_193_ ), .A4(\EXU/ALU/_194_ ), .ZN(\EXU/ALU/_195_ ) );
NAND4_X1 \EXU/ALU/_488_ ( .A1(\EXU/ALU/_186_ ), .A2(fanout_net_12 ), .A3(fanout_net_13 ), .A4(\EXU/ALU/_146_ ), .ZN(\EXU/ALU/_196_ ) );
AND2_X1 \EXU/ALU/_489_ ( .A1(\EXU/ALU/_195_ ), .A2(\EXU/ALU/_196_ ), .ZN(\EXU/ALU/_197_ ) );
BUF_X4 \EXU/ALU/_490_ ( .A(\EXU/ALU/_193_ ), .Z(\EXU/ALU/_198_ ) );
BUF_X4 \EXU/ALU/_491_ ( .A(\EXU/ALU/_174_ ), .Z(\EXU/ALU/_199_ ) );
NAND3_X1 \EXU/ALU/_492_ ( .A1(\EXU/ALU/_198_ ), .A2(\EXU/ALU/_199_ ), .A3(\EXU/ALU/_013_ ), .ZN(\EXU/ALU/_200_ ) );
AOI22_X1 \EXU/ALU/_493_ ( .A1(\EXU/ALU/_183_ ), .A2(\EXU/ALU/_192_ ), .B1(\EXU/ALU/_050_ ), .B2(\EXU/ALU/_190_ ), .ZN(\EXU/ALU/_201_ ) );
BUF_X4 \EXU/ALU/_494_ ( .A(\EXU/ALU/_185_ ), .Z(\EXU/ALU/_202_ ) );
NAND4_X1 \EXU/ALU/_495_ ( .A1(\EXU/ALU/_202_ ), .A2(fanout_net_14 ), .A3(\EXU/ALU/_146_ ), .A4(\EXU/ALU/_114_ ), .ZN(\EXU/ALU/_203_ ) );
NAND4_X1 \EXU/ALU/_496_ ( .A1(\EXU/ALU/_197_ ), .A2(\EXU/ALU/_200_ ), .A3(\EXU/ALU/_201_ ), .A4(\EXU/ALU/_203_ ), .ZN(\EXU/ALU/_082_ ) );
OR2_X1 \EXU/ALU/_497_ ( .A1(\EXU/ALU/_157_ ), .A2(\EXU/ALU/_125_ ), .ZN(\EXU/ALU/_204_ ) );
NAND2_X1 \EXU/ALU/_498_ ( .A1(\EXU/ALU/_157_ ), .A2(\EXU/ALU/_125_ ), .ZN(\EXU/ALU/_205_ ) );
NAND4_X1 \EXU/ALU/_499_ ( .A1(\EXU/ALU/_204_ ), .A2(fanout_net_14 ), .A3(\EXU/ALU/_193_ ), .A4(\EXU/ALU/_205_ ), .ZN(\EXU/ALU/_206_ ) );
NAND4_X1 \EXU/ALU/_500_ ( .A1(\EXU/ALU/_186_ ), .A2(fanout_net_12 ), .A3(fanout_net_13 ), .A4(\EXU/ALU/_157_ ), .ZN(\EXU/ALU/_207_ ) );
AND2_X1 \EXU/ALU/_501_ ( .A1(\EXU/ALU/_206_ ), .A2(\EXU/ALU/_207_ ), .ZN(\EXU/ALU/_208_ ) );
NAND3_X1 \EXU/ALU/_502_ ( .A1(\EXU/ALU/_198_ ), .A2(\EXU/ALU/_199_ ), .A3(\EXU/ALU/_024_ ), .ZN(\EXU/ALU/_209_ ) );
AOI22_X2 \EXU/ALU/_503_ ( .A1(\EXU/ALU/_183_ ), .A2(\EXU/ALU/_204_ ), .B1(\EXU/ALU/_061_ ), .B2(\EXU/ALU/_190_ ), .ZN(\EXU/ALU/_210_ ) );
NAND4_X1 \EXU/ALU/_504_ ( .A1(\EXU/ALU/_202_ ), .A2(fanout_net_14 ), .A3(\EXU/ALU/_157_ ), .A4(\EXU/ALU/_125_ ), .ZN(\EXU/ALU/_211_ ) );
NAND4_X1 \EXU/ALU/_505_ ( .A1(\EXU/ALU/_208_ ), .A2(\EXU/ALU/_209_ ), .A3(\EXU/ALU/_210_ ), .A4(\EXU/ALU/_211_ ), .ZN(\EXU/ALU/_093_ ) );
OR2_X1 \EXU/ALU/_506_ ( .A1(\EXU/ALU/_160_ ), .A2(\EXU/ALU/_128_ ), .ZN(\EXU/ALU/_212_ ) );
NAND2_X1 \EXU/ALU/_507_ ( .A1(\EXU/ALU/_160_ ), .A2(\EXU/ALU/_128_ ), .ZN(\EXU/ALU/_213_ ) );
NAND4_X1 \EXU/ALU/_508_ ( .A1(\EXU/ALU/_212_ ), .A2(fanout_net_14 ), .A3(\EXU/ALU/_193_ ), .A4(\EXU/ALU/_213_ ), .ZN(\EXU/ALU/_214_ ) );
NAND4_X1 \EXU/ALU/_509_ ( .A1(\EXU/ALU/_186_ ), .A2(fanout_net_12 ), .A3(fanout_net_13 ), .A4(\EXU/ALU/_160_ ), .ZN(\EXU/ALU/_215_ ) );
AND2_X1 \EXU/ALU/_510_ ( .A1(\EXU/ALU/_214_ ), .A2(\EXU/ALU/_215_ ), .ZN(\EXU/ALU/_216_ ) );
NAND3_X1 \EXU/ALU/_511_ ( .A1(\EXU/ALU/_198_ ), .A2(\EXU/ALU/_199_ ), .A3(\EXU/ALU/_027_ ), .ZN(\EXU/ALU/_217_ ) );
AOI22_X2 \EXU/ALU/_512_ ( .A1(\EXU/ALU/_183_ ), .A2(\EXU/ALU/_212_ ), .B1(\EXU/ALU/_064_ ), .B2(\EXU/ALU/_190_ ), .ZN(\EXU/ALU/_218_ ) );
NAND4_X1 \EXU/ALU/_513_ ( .A1(\EXU/ALU/_202_ ), .A2(fanout_net_14 ), .A3(\EXU/ALU/_160_ ), .A4(\EXU/ALU/_128_ ), .ZN(\EXU/ALU/_219_ ) );
NAND4_X1 \EXU/ALU/_514_ ( .A1(\EXU/ALU/_216_ ), .A2(\EXU/ALU/_217_ ), .A3(\EXU/ALU/_218_ ), .A4(\EXU/ALU/_219_ ), .ZN(\EXU/ALU/_096_ ) );
OR2_X1 \EXU/ALU/_515_ ( .A1(\EXU/ALU/_161_ ), .A2(\EXU/ALU/_129_ ), .ZN(\EXU/ALU/_220_ ) );
NAND2_X1 \EXU/ALU/_516_ ( .A1(\EXU/ALU/_161_ ), .A2(\EXU/ALU/_129_ ), .ZN(\EXU/ALU/_221_ ) );
NAND4_X1 \EXU/ALU/_517_ ( .A1(\EXU/ALU/_220_ ), .A2(fanout_net_14 ), .A3(\EXU/ALU/_193_ ), .A4(\EXU/ALU/_221_ ), .ZN(\EXU/ALU/_222_ ) );
NAND4_X1 \EXU/ALU/_518_ ( .A1(\EXU/ALU/_186_ ), .A2(fanout_net_12 ), .A3(fanout_net_13 ), .A4(\EXU/ALU/_161_ ), .ZN(\EXU/ALU/_223_ ) );
AND2_X1 \EXU/ALU/_519_ ( .A1(\EXU/ALU/_222_ ), .A2(\EXU/ALU/_223_ ), .ZN(\EXU/ALU/_224_ ) );
NAND3_X1 \EXU/ALU/_520_ ( .A1(\EXU/ALU/_198_ ), .A2(\EXU/ALU/_199_ ), .A3(\EXU/ALU/_028_ ), .ZN(\EXU/ALU/_225_ ) );
AOI22_X1 \EXU/ALU/_521_ ( .A1(\EXU/ALU/_183_ ), .A2(\EXU/ALU/_220_ ), .B1(\EXU/ALU/_065_ ), .B2(\EXU/ALU/_190_ ), .ZN(\EXU/ALU/_226_ ) );
NAND4_X1 \EXU/ALU/_522_ ( .A1(\EXU/ALU/_202_ ), .A2(fanout_net_14 ), .A3(\EXU/ALU/_161_ ), .A4(\EXU/ALU/_129_ ), .ZN(\EXU/ALU/_227_ ) );
NAND4_X1 \EXU/ALU/_523_ ( .A1(\EXU/ALU/_224_ ), .A2(\EXU/ALU/_225_ ), .A3(\EXU/ALU/_226_ ), .A4(\EXU/ALU/_227_ ), .ZN(\EXU/ALU/_097_ ) );
OR2_X1 \EXU/ALU/_524_ ( .A1(\EXU/ALU/_162_ ), .A2(\EXU/ALU/_130_ ), .ZN(\EXU/ALU/_228_ ) );
NAND2_X1 \EXU/ALU/_525_ ( .A1(\EXU/ALU/_162_ ), .A2(\EXU/ALU/_130_ ), .ZN(\EXU/ALU/_229_ ) );
NAND4_X1 \EXU/ALU/_526_ ( .A1(\EXU/ALU/_228_ ), .A2(fanout_net_14 ), .A3(\EXU/ALU/_193_ ), .A4(\EXU/ALU/_229_ ), .ZN(\EXU/ALU/_230_ ) );
NAND4_X1 \EXU/ALU/_527_ ( .A1(\EXU/ALU/_186_ ), .A2(fanout_net_12 ), .A3(fanout_net_13 ), .A4(\EXU/ALU/_162_ ), .ZN(\EXU/ALU/_231_ ) );
AND2_X1 \EXU/ALU/_528_ ( .A1(\EXU/ALU/_230_ ), .A2(\EXU/ALU/_231_ ), .ZN(\EXU/ALU/_232_ ) );
NAND3_X1 \EXU/ALU/_529_ ( .A1(\EXU/ALU/_198_ ), .A2(\EXU/ALU/_199_ ), .A3(\EXU/ALU/_029_ ), .ZN(\EXU/ALU/_233_ ) );
AOI22_X1 \EXU/ALU/_530_ ( .A1(\EXU/ALU/_183_ ), .A2(\EXU/ALU/_228_ ), .B1(\EXU/ALU/_066_ ), .B2(\EXU/ALU/_190_ ), .ZN(\EXU/ALU/_234_ ) );
NAND4_X1 \EXU/ALU/_531_ ( .A1(\EXU/ALU/_202_ ), .A2(fanout_net_14 ), .A3(\EXU/ALU/_162_ ), .A4(\EXU/ALU/_130_ ), .ZN(\EXU/ALU/_235_ ) );
NAND4_X1 \EXU/ALU/_532_ ( .A1(\EXU/ALU/_232_ ), .A2(\EXU/ALU/_233_ ), .A3(\EXU/ALU/_234_ ), .A4(\EXU/ALU/_235_ ), .ZN(\EXU/ALU/_098_ ) );
OR2_X1 \EXU/ALU/_533_ ( .A1(\EXU/ALU/_163_ ), .A2(\EXU/ALU/_131_ ), .ZN(\EXU/ALU/_236_ ) );
NAND2_X1 \EXU/ALU/_534_ ( .A1(\EXU/ALU/_163_ ), .A2(\EXU/ALU/_131_ ), .ZN(\EXU/ALU/_237_ ) );
NAND4_X1 \EXU/ALU/_535_ ( .A1(\EXU/ALU/_236_ ), .A2(fanout_net_14 ), .A3(\EXU/ALU/_193_ ), .A4(\EXU/ALU/_237_ ), .ZN(\EXU/ALU/_238_ ) );
NAND4_X1 \EXU/ALU/_536_ ( .A1(\EXU/ALU/_186_ ), .A2(fanout_net_12 ), .A3(fanout_net_13 ), .A4(\EXU/ALU/_163_ ), .ZN(\EXU/ALU/_239_ ) );
AND2_X1 \EXU/ALU/_537_ ( .A1(\EXU/ALU/_238_ ), .A2(\EXU/ALU/_239_ ), .ZN(\EXU/ALU/_240_ ) );
NAND3_X1 \EXU/ALU/_538_ ( .A1(\EXU/ALU/_198_ ), .A2(\EXU/ALU/_199_ ), .A3(\EXU/ALU/_030_ ), .ZN(\EXU/ALU/_241_ ) );
AOI22_X2 \EXU/ALU/_539_ ( .A1(\EXU/ALU/_183_ ), .A2(\EXU/ALU/_236_ ), .B1(\EXU/ALU/_067_ ), .B2(\EXU/ALU/_190_ ), .ZN(\EXU/ALU/_242_ ) );
NAND4_X1 \EXU/ALU/_540_ ( .A1(\EXU/ALU/_202_ ), .A2(fanout_net_14 ), .A3(\EXU/ALU/_163_ ), .A4(\EXU/ALU/_131_ ), .ZN(\EXU/ALU/_243_ ) );
NAND4_X1 \EXU/ALU/_541_ ( .A1(\EXU/ALU/_240_ ), .A2(\EXU/ALU/_241_ ), .A3(\EXU/ALU/_242_ ), .A4(\EXU/ALU/_243_ ), .ZN(\EXU/ALU/_099_ ) );
OR2_X1 \EXU/ALU/_542_ ( .A1(\EXU/ALU/_164_ ), .A2(\EXU/ALU/_132_ ), .ZN(\EXU/ALU/_244_ ) );
BUF_X4 \EXU/ALU/_543_ ( .A(\EXU/ALU/_178_ ), .Z(\EXU/ALU/_245_ ) );
NAND2_X1 \EXU/ALU/_544_ ( .A1(\EXU/ALU/_164_ ), .A2(\EXU/ALU/_132_ ), .ZN(\EXU/ALU/_246_ ) );
NAND4_X1 \EXU/ALU/_545_ ( .A1(\EXU/ALU/_244_ ), .A2(fanout_net_14 ), .A3(\EXU/ALU/_245_ ), .A4(\EXU/ALU/_246_ ), .ZN(\EXU/ALU/_247_ ) );
NAND4_X1 \EXU/ALU/_546_ ( .A1(\EXU/ALU/_186_ ), .A2(fanout_net_12 ), .A3(fanout_net_13 ), .A4(\EXU/ALU/_164_ ), .ZN(\EXU/ALU/_248_ ) );
AND2_X1 \EXU/ALU/_547_ ( .A1(\EXU/ALU/_247_ ), .A2(\EXU/ALU/_248_ ), .ZN(\EXU/ALU/_249_ ) );
NAND3_X1 \EXU/ALU/_548_ ( .A1(\EXU/ALU/_198_ ), .A2(\EXU/ALU/_199_ ), .A3(\EXU/ALU/_031_ ), .ZN(\EXU/ALU/_250_ ) );
AOI22_X2 \EXU/ALU/_549_ ( .A1(\EXU/ALU/_183_ ), .A2(\EXU/ALU/_244_ ), .B1(\EXU/ALU/_068_ ), .B2(\EXU/ALU/_190_ ), .ZN(\EXU/ALU/_251_ ) );
NAND4_X1 \EXU/ALU/_550_ ( .A1(\EXU/ALU/_202_ ), .A2(fanout_net_14 ), .A3(\EXU/ALU/_164_ ), .A4(\EXU/ALU/_132_ ), .ZN(\EXU/ALU/_252_ ) );
NAND4_X1 \EXU/ALU/_551_ ( .A1(\EXU/ALU/_249_ ), .A2(\EXU/ALU/_250_ ), .A3(\EXU/ALU/_251_ ), .A4(\EXU/ALU/_252_ ), .ZN(\EXU/ALU/_100_ ) );
OR2_X1 \EXU/ALU/_552_ ( .A1(\EXU/ALU/_165_ ), .A2(\EXU/ALU/_133_ ), .ZN(\EXU/ALU/_253_ ) );
NAND2_X1 \EXU/ALU/_553_ ( .A1(\EXU/ALU/_165_ ), .A2(\EXU/ALU/_133_ ), .ZN(\EXU/ALU/_254_ ) );
NAND4_X1 \EXU/ALU/_554_ ( .A1(\EXU/ALU/_253_ ), .A2(fanout_net_14 ), .A3(\EXU/ALU/_245_ ), .A4(\EXU/ALU/_254_ ), .ZN(\EXU/ALU/_255_ ) );
NAND4_X1 \EXU/ALU/_555_ ( .A1(\EXU/ALU/_186_ ), .A2(fanout_net_12 ), .A3(fanout_net_13 ), .A4(\EXU/ALU/_165_ ), .ZN(\EXU/ALU/_256_ ) );
AND2_X1 \EXU/ALU/_556_ ( .A1(\EXU/ALU/_255_ ), .A2(\EXU/ALU/_256_ ), .ZN(\EXU/ALU/_257_ ) );
NAND3_X1 \EXU/ALU/_557_ ( .A1(\EXU/ALU/_198_ ), .A2(\EXU/ALU/_199_ ), .A3(\EXU/ALU/_032_ ), .ZN(\EXU/ALU/_258_ ) );
AOI22_X1 \EXU/ALU/_558_ ( .A1(\EXU/ALU/_183_ ), .A2(\EXU/ALU/_253_ ), .B1(\EXU/ALU/_069_ ), .B2(\EXU/ALU/_190_ ), .ZN(\EXU/ALU/_259_ ) );
NAND4_X1 \EXU/ALU/_559_ ( .A1(\EXU/ALU/_202_ ), .A2(fanout_net_14 ), .A3(\EXU/ALU/_165_ ), .A4(\EXU/ALU/_133_ ), .ZN(\EXU/ALU/_260_ ) );
NAND4_X1 \EXU/ALU/_560_ ( .A1(\EXU/ALU/_257_ ), .A2(\EXU/ALU/_258_ ), .A3(\EXU/ALU/_259_ ), .A4(\EXU/ALU/_260_ ), .ZN(\EXU/ALU/_101_ ) );
OR2_X1 \EXU/ALU/_561_ ( .A1(\EXU/ALU/_166_ ), .A2(\EXU/ALU/_134_ ), .ZN(\EXU/ALU/_261_ ) );
NAND2_X1 \EXU/ALU/_562_ ( .A1(\EXU/ALU/_166_ ), .A2(\EXU/ALU/_134_ ), .ZN(\EXU/ALU/_262_ ) );
NAND4_X1 \EXU/ALU/_563_ ( .A1(\EXU/ALU/_261_ ), .A2(fanout_net_14 ), .A3(\EXU/ALU/_245_ ), .A4(\EXU/ALU/_262_ ), .ZN(\EXU/ALU/_263_ ) );
BUF_X8 \EXU/ALU/_564_ ( .A(\EXU/ALU/_174_ ), .Z(\EXU/ALU/_264_ ) );
NAND4_X1 \EXU/ALU/_565_ ( .A1(\EXU/ALU/_264_ ), .A2(fanout_net_12 ), .A3(fanout_net_13 ), .A4(\EXU/ALU/_166_ ), .ZN(\EXU/ALU/_265_ ) );
AND2_X1 \EXU/ALU/_566_ ( .A1(\EXU/ALU/_263_ ), .A2(\EXU/ALU/_265_ ), .ZN(\EXU/ALU/_266_ ) );
NAND3_X1 \EXU/ALU/_567_ ( .A1(\EXU/ALU/_198_ ), .A2(\EXU/ALU/_199_ ), .A3(\EXU/ALU/_033_ ), .ZN(\EXU/ALU/_267_ ) );
AOI22_X1 \EXU/ALU/_568_ ( .A1(\EXU/ALU/_183_ ), .A2(\EXU/ALU/_261_ ), .B1(\EXU/ALU/_070_ ), .B2(\EXU/ALU/_190_ ), .ZN(\EXU/ALU/_268_ ) );
NAND4_X1 \EXU/ALU/_569_ ( .A1(\EXU/ALU/_202_ ), .A2(fanout_net_14 ), .A3(\EXU/ALU/_166_ ), .A4(\EXU/ALU/_134_ ), .ZN(\EXU/ALU/_269_ ) );
NAND4_X1 \EXU/ALU/_570_ ( .A1(\EXU/ALU/_266_ ), .A2(\EXU/ALU/_267_ ), .A3(\EXU/ALU/_268_ ), .A4(\EXU/ALU/_269_ ), .ZN(\EXU/ALU/_102_ ) );
OR2_X1 \EXU/ALU/_571_ ( .A1(\EXU/ALU/_136_ ), .A2(\EXU/ALU/_104_ ), .ZN(\EXU/ALU/_270_ ) );
NAND2_X1 \EXU/ALU/_572_ ( .A1(\EXU/ALU/_136_ ), .A2(\EXU/ALU/_104_ ), .ZN(\EXU/ALU/_271_ ) );
NAND4_X1 \EXU/ALU/_573_ ( .A1(\EXU/ALU/_270_ ), .A2(fanout_net_14 ), .A3(\EXU/ALU/_245_ ), .A4(\EXU/ALU/_271_ ), .ZN(\EXU/ALU/_272_ ) );
NAND4_X1 \EXU/ALU/_574_ ( .A1(\EXU/ALU/_264_ ), .A2(fanout_net_12 ), .A3(fanout_net_13 ), .A4(\EXU/ALU/_136_ ), .ZN(\EXU/ALU/_273_ ) );
AND2_X1 \EXU/ALU/_575_ ( .A1(\EXU/ALU/_272_ ), .A2(\EXU/ALU/_273_ ), .ZN(\EXU/ALU/_274_ ) );
NAND3_X1 \EXU/ALU/_576_ ( .A1(\EXU/ALU/_198_ ), .A2(\EXU/ALU/_199_ ), .A3(\EXU/ALU/_003_ ), .ZN(\EXU/ALU/_275_ ) );
BUF_X4 \EXU/ALU/_577_ ( .A(\EXU/ALU/_182_ ), .Z(\EXU/ALU/_276_ ) );
BUF_X4 \EXU/ALU/_578_ ( .A(\EXU/ALU/_189_ ), .Z(\EXU/ALU/_277_ ) );
AOI22_X1 \EXU/ALU/_579_ ( .A1(\EXU/ALU/_276_ ), .A2(\EXU/ALU/_270_ ), .B1(\EXU/ALU/_040_ ), .B2(\EXU/ALU/_277_ ), .ZN(\EXU/ALU/_278_ ) );
NAND4_X1 \EXU/ALU/_580_ ( .A1(\EXU/ALU/_202_ ), .A2(fanout_net_14 ), .A3(\EXU/ALU/_136_ ), .A4(\EXU/ALU/_104_ ), .ZN(\EXU/ALU/_279_ ) );
NAND4_X1 \EXU/ALU/_581_ ( .A1(\EXU/ALU/_274_ ), .A2(\EXU/ALU/_275_ ), .A3(\EXU/ALU/_278_ ), .A4(\EXU/ALU/_279_ ), .ZN(\EXU/ALU/_072_ ) );
OR2_X1 \EXU/ALU/_582_ ( .A1(\EXU/ALU/_137_ ), .A2(\EXU/ALU/_105_ ), .ZN(\EXU/ALU/_280_ ) );
NAND2_X1 \EXU/ALU/_583_ ( .A1(\EXU/ALU/_137_ ), .A2(\EXU/ALU/_105_ ), .ZN(\EXU/ALU/_281_ ) );
NAND4_X1 \EXU/ALU/_584_ ( .A1(\EXU/ALU/_280_ ), .A2(fanout_net_14 ), .A3(\EXU/ALU/_245_ ), .A4(\EXU/ALU/_281_ ), .ZN(\EXU/ALU/_282_ ) );
NAND4_X1 \EXU/ALU/_585_ ( .A1(\EXU/ALU/_264_ ), .A2(fanout_net_12 ), .A3(fanout_net_13 ), .A4(\EXU/ALU/_137_ ), .ZN(\EXU/ALU/_283_ ) );
AND2_X1 \EXU/ALU/_586_ ( .A1(\EXU/ALU/_282_ ), .A2(\EXU/ALU/_283_ ), .ZN(\EXU/ALU/_284_ ) );
BUF_X4 \EXU/ALU/_587_ ( .A(\EXU/ALU/_193_ ), .Z(\EXU/ALU/_285_ ) );
BUF_X4 \EXU/ALU/_588_ ( .A(\EXU/ALU/_174_ ), .Z(\EXU/ALU/_286_ ) );
NAND3_X1 \EXU/ALU/_589_ ( .A1(\EXU/ALU/_285_ ), .A2(\EXU/ALU/_286_ ), .A3(\EXU/ALU/_004_ ), .ZN(\EXU/ALU/_287_ ) );
AOI22_X1 \EXU/ALU/_590_ ( .A1(\EXU/ALU/_276_ ), .A2(\EXU/ALU/_280_ ), .B1(\EXU/ALU/_041_ ), .B2(\EXU/ALU/_277_ ), .ZN(\EXU/ALU/_288_ ) );
BUF_X4 \EXU/ALU/_591_ ( .A(\EXU/ALU/_185_ ), .Z(\EXU/ALU/_289_ ) );
NAND4_X1 \EXU/ALU/_592_ ( .A1(\EXU/ALU/_289_ ), .A2(fanout_net_14 ), .A3(\EXU/ALU/_137_ ), .A4(\EXU/ALU/_105_ ), .ZN(\EXU/ALU/_290_ ) );
NAND4_X1 \EXU/ALU/_593_ ( .A1(\EXU/ALU/_284_ ), .A2(\EXU/ALU/_287_ ), .A3(\EXU/ALU/_288_ ), .A4(\EXU/ALU/_290_ ), .ZN(\EXU/ALU/_073_ ) );
OR2_X1 \EXU/ALU/_594_ ( .A1(\EXU/ALU/_138_ ), .A2(\EXU/ALU/_106_ ), .ZN(\EXU/ALU/_291_ ) );
NAND2_X1 \EXU/ALU/_595_ ( .A1(\EXU/ALU/_138_ ), .A2(\EXU/ALU/_106_ ), .ZN(\EXU/ALU/_292_ ) );
NAND4_X1 \EXU/ALU/_596_ ( .A1(\EXU/ALU/_291_ ), .A2(fanout_net_14 ), .A3(\EXU/ALU/_245_ ), .A4(\EXU/ALU/_292_ ), .ZN(\EXU/ALU/_293_ ) );
NAND4_X1 \EXU/ALU/_597_ ( .A1(\EXU/ALU/_264_ ), .A2(fanout_net_12 ), .A3(fanout_net_13 ), .A4(\EXU/ALU/_138_ ), .ZN(\EXU/ALU/_294_ ) );
AND2_X1 \EXU/ALU/_598_ ( .A1(\EXU/ALU/_293_ ), .A2(\EXU/ALU/_294_ ), .ZN(\EXU/ALU/_295_ ) );
NAND3_X1 \EXU/ALU/_599_ ( .A1(\EXU/ALU/_285_ ), .A2(\EXU/ALU/_286_ ), .A3(\EXU/ALU/_005_ ), .ZN(\EXU/ALU/_296_ ) );
AOI22_X1 \EXU/ALU/_600_ ( .A1(\EXU/ALU/_276_ ), .A2(\EXU/ALU/_291_ ), .B1(\EXU/ALU/_042_ ), .B2(\EXU/ALU/_277_ ), .ZN(\EXU/ALU/_297_ ) );
NAND4_X1 \EXU/ALU/_601_ ( .A1(\EXU/ALU/_289_ ), .A2(fanout_net_14 ), .A3(\EXU/ALU/_138_ ), .A4(\EXU/ALU/_106_ ), .ZN(\EXU/ALU/_298_ ) );
NAND4_X1 \EXU/ALU/_602_ ( .A1(\EXU/ALU/_295_ ), .A2(\EXU/ALU/_296_ ), .A3(\EXU/ALU/_297_ ), .A4(\EXU/ALU/_298_ ), .ZN(\EXU/ALU/_074_ ) );
OR2_X1 \EXU/ALU/_603_ ( .A1(\EXU/ALU/_139_ ), .A2(\EXU/ALU/_107_ ), .ZN(\EXU/ALU/_299_ ) );
NAND2_X1 \EXU/ALU/_604_ ( .A1(\EXU/ALU/_139_ ), .A2(\EXU/ALU/_107_ ), .ZN(\EXU/ALU/_300_ ) );
NAND4_X1 \EXU/ALU/_605_ ( .A1(\EXU/ALU/_299_ ), .A2(fanout_net_14 ), .A3(\EXU/ALU/_245_ ), .A4(\EXU/ALU/_300_ ), .ZN(\EXU/ALU/_301_ ) );
NAND4_X1 \EXU/ALU/_606_ ( .A1(\EXU/ALU/_264_ ), .A2(fanout_net_12 ), .A3(fanout_net_13 ), .A4(\EXU/ALU/_139_ ), .ZN(\EXU/ALU/_302_ ) );
AND2_X1 \EXU/ALU/_607_ ( .A1(\EXU/ALU/_301_ ), .A2(\EXU/ALU/_302_ ), .ZN(\EXU/ALU/_303_ ) );
NAND3_X1 \EXU/ALU/_608_ ( .A1(\EXU/ALU/_285_ ), .A2(\EXU/ALU/_286_ ), .A3(\EXU/ALU/_006_ ), .ZN(\EXU/ALU/_304_ ) );
AOI22_X1 \EXU/ALU/_609_ ( .A1(\EXU/ALU/_276_ ), .A2(\EXU/ALU/_299_ ), .B1(\EXU/ALU/_043_ ), .B2(\EXU/ALU/_277_ ), .ZN(\EXU/ALU/_305_ ) );
NAND4_X1 \EXU/ALU/_610_ ( .A1(\EXU/ALU/_289_ ), .A2(fanout_net_14 ), .A3(\EXU/ALU/_139_ ), .A4(\EXU/ALU/_107_ ), .ZN(\EXU/ALU/_306_ ) );
NAND4_X1 \EXU/ALU/_611_ ( .A1(\EXU/ALU/_303_ ), .A2(\EXU/ALU/_304_ ), .A3(\EXU/ALU/_305_ ), .A4(\EXU/ALU/_306_ ), .ZN(\EXU/ALU/_075_ ) );
OR2_X1 \EXU/ALU/_612_ ( .A1(\EXU/ALU/_140_ ), .A2(\EXU/ALU/_108_ ), .ZN(\EXU/ALU/_307_ ) );
NAND2_X1 \EXU/ALU/_613_ ( .A1(\EXU/ALU/_140_ ), .A2(\EXU/ALU/_108_ ), .ZN(\EXU/ALU/_308_ ) );
NAND4_X1 \EXU/ALU/_614_ ( .A1(\EXU/ALU/_307_ ), .A2(fanout_net_14 ), .A3(\EXU/ALU/_245_ ), .A4(\EXU/ALU/_308_ ), .ZN(\EXU/ALU/_309_ ) );
NAND4_X1 \EXU/ALU/_615_ ( .A1(\EXU/ALU/_264_ ), .A2(fanout_net_12 ), .A3(fanout_net_13 ), .A4(\EXU/ALU/_140_ ), .ZN(\EXU/ALU/_310_ ) );
AND2_X1 \EXU/ALU/_616_ ( .A1(\EXU/ALU/_309_ ), .A2(\EXU/ALU/_310_ ), .ZN(\EXU/ALU/_311_ ) );
NAND3_X1 \EXU/ALU/_617_ ( .A1(\EXU/ALU/_285_ ), .A2(\EXU/ALU/_286_ ), .A3(\EXU/ALU/_007_ ), .ZN(\EXU/ALU/_312_ ) );
AOI22_X1 \EXU/ALU/_618_ ( .A1(\EXU/ALU/_276_ ), .A2(\EXU/ALU/_307_ ), .B1(\EXU/ALU/_044_ ), .B2(\EXU/ALU/_277_ ), .ZN(\EXU/ALU/_313_ ) );
NAND4_X1 \EXU/ALU/_619_ ( .A1(\EXU/ALU/_289_ ), .A2(fanout_net_14 ), .A3(\EXU/ALU/_140_ ), .A4(\EXU/ALU/_108_ ), .ZN(\EXU/ALU/_314_ ) );
NAND4_X1 \EXU/ALU/_620_ ( .A1(\EXU/ALU/_311_ ), .A2(\EXU/ALU/_312_ ), .A3(\EXU/ALU/_313_ ), .A4(\EXU/ALU/_314_ ), .ZN(\EXU/ALU/_076_ ) );
OR2_X1 \EXU/ALU/_621_ ( .A1(\EXU/ALU/_141_ ), .A2(\EXU/ALU/_109_ ), .ZN(\EXU/ALU/_315_ ) );
NAND2_X1 \EXU/ALU/_622_ ( .A1(\EXU/ALU/_141_ ), .A2(\EXU/ALU/_109_ ), .ZN(\EXU/ALU/_316_ ) );
NAND4_X1 \EXU/ALU/_623_ ( .A1(\EXU/ALU/_315_ ), .A2(fanout_net_15 ), .A3(\EXU/ALU/_245_ ), .A4(\EXU/ALU/_316_ ), .ZN(\EXU/ALU/_317_ ) );
NAND4_X1 \EXU/ALU/_624_ ( .A1(\EXU/ALU/_264_ ), .A2(fanout_net_12 ), .A3(fanout_net_13 ), .A4(\EXU/ALU/_141_ ), .ZN(\EXU/ALU/_318_ ) );
AND2_X1 \EXU/ALU/_625_ ( .A1(\EXU/ALU/_317_ ), .A2(\EXU/ALU/_318_ ), .ZN(\EXU/ALU/_319_ ) );
NAND3_X1 \EXU/ALU/_626_ ( .A1(\EXU/ALU/_285_ ), .A2(\EXU/ALU/_286_ ), .A3(\EXU/ALU/_008_ ), .ZN(\EXU/ALU/_320_ ) );
AOI22_X1 \EXU/ALU/_627_ ( .A1(\EXU/ALU/_276_ ), .A2(\EXU/ALU/_315_ ), .B1(\EXU/ALU/_045_ ), .B2(\EXU/ALU/_277_ ), .ZN(\EXU/ALU/_321_ ) );
NAND4_X1 \EXU/ALU/_628_ ( .A1(\EXU/ALU/_289_ ), .A2(fanout_net_15 ), .A3(\EXU/ALU/_141_ ), .A4(\EXU/ALU/_109_ ), .ZN(\EXU/ALU/_322_ ) );
NAND4_X1 \EXU/ALU/_629_ ( .A1(\EXU/ALU/_319_ ), .A2(\EXU/ALU/_320_ ), .A3(\EXU/ALU/_321_ ), .A4(\EXU/ALU/_322_ ), .ZN(\EXU/ALU/_077_ ) );
OR2_X1 \EXU/ALU/_630_ ( .A1(\EXU/ALU/_142_ ), .A2(\EXU/ALU/_110_ ), .ZN(\EXU/ALU/_323_ ) );
NAND2_X1 \EXU/ALU/_631_ ( .A1(\EXU/ALU/_142_ ), .A2(\EXU/ALU/_110_ ), .ZN(\EXU/ALU/_324_ ) );
NAND4_X1 \EXU/ALU/_632_ ( .A1(\EXU/ALU/_323_ ), .A2(fanout_net_15 ), .A3(\EXU/ALU/_245_ ), .A4(\EXU/ALU/_324_ ), .ZN(\EXU/ALU/_325_ ) );
NAND4_X1 \EXU/ALU/_633_ ( .A1(\EXU/ALU/_264_ ), .A2(fanout_net_12 ), .A3(fanout_net_13 ), .A4(\EXU/ALU/_142_ ), .ZN(\EXU/ALU/_326_ ) );
AND2_X1 \EXU/ALU/_634_ ( .A1(\EXU/ALU/_325_ ), .A2(\EXU/ALU/_326_ ), .ZN(\EXU/ALU/_327_ ) );
NAND3_X1 \EXU/ALU/_635_ ( .A1(\EXU/ALU/_285_ ), .A2(\EXU/ALU/_286_ ), .A3(\EXU/ALU/_009_ ), .ZN(\EXU/ALU/_328_ ) );
AOI22_X1 \EXU/ALU/_636_ ( .A1(\EXU/ALU/_276_ ), .A2(\EXU/ALU/_323_ ), .B1(\EXU/ALU/_046_ ), .B2(\EXU/ALU/_277_ ), .ZN(\EXU/ALU/_329_ ) );
NAND4_X1 \EXU/ALU/_637_ ( .A1(\EXU/ALU/_289_ ), .A2(fanout_net_15 ), .A3(\EXU/ALU/_142_ ), .A4(\EXU/ALU/_110_ ), .ZN(\EXU/ALU/_330_ ) );
NAND4_X1 \EXU/ALU/_638_ ( .A1(\EXU/ALU/_327_ ), .A2(\EXU/ALU/_328_ ), .A3(\EXU/ALU/_329_ ), .A4(\EXU/ALU/_330_ ), .ZN(\EXU/ALU/_078_ ) );
OR2_X1 \EXU/ALU/_639_ ( .A1(\EXU/ALU/_143_ ), .A2(\EXU/ALU/_111_ ), .ZN(\EXU/ALU/_331_ ) );
BUF_X4 \EXU/ALU/_640_ ( .A(\EXU/ALU/_178_ ), .Z(\EXU/ALU/_332_ ) );
NAND2_X1 \EXU/ALU/_641_ ( .A1(\EXU/ALU/_143_ ), .A2(\EXU/ALU/_111_ ), .ZN(\EXU/ALU/_333_ ) );
NAND4_X1 \EXU/ALU/_642_ ( .A1(\EXU/ALU/_331_ ), .A2(fanout_net_15 ), .A3(\EXU/ALU/_332_ ), .A4(\EXU/ALU/_333_ ), .ZN(\EXU/ALU/_334_ ) );
NAND4_X1 \EXU/ALU/_643_ ( .A1(\EXU/ALU/_264_ ), .A2(fanout_net_12 ), .A3(fanout_net_13 ), .A4(\EXU/ALU/_143_ ), .ZN(\EXU/ALU/_335_ ) );
AND2_X1 \EXU/ALU/_644_ ( .A1(\EXU/ALU/_334_ ), .A2(\EXU/ALU/_335_ ), .ZN(\EXU/ALU/_336_ ) );
NAND3_X1 \EXU/ALU/_645_ ( .A1(\EXU/ALU/_285_ ), .A2(\EXU/ALU/_286_ ), .A3(\EXU/ALU/_010_ ), .ZN(\EXU/ALU/_337_ ) );
AOI22_X1 \EXU/ALU/_646_ ( .A1(\EXU/ALU/_276_ ), .A2(\EXU/ALU/_331_ ), .B1(\EXU/ALU/_047_ ), .B2(\EXU/ALU/_277_ ), .ZN(\EXU/ALU/_338_ ) );
NAND4_X1 \EXU/ALU/_647_ ( .A1(\EXU/ALU/_289_ ), .A2(fanout_net_15 ), .A3(\EXU/ALU/_143_ ), .A4(\EXU/ALU/_111_ ), .ZN(\EXU/ALU/_339_ ) );
NAND4_X1 \EXU/ALU/_648_ ( .A1(\EXU/ALU/_336_ ), .A2(\EXU/ALU/_337_ ), .A3(\EXU/ALU/_338_ ), .A4(\EXU/ALU/_339_ ), .ZN(\EXU/ALU/_079_ ) );
OR2_X1 \EXU/ALU/_649_ ( .A1(\EXU/ALU/_144_ ), .A2(\EXU/ALU/_112_ ), .ZN(\EXU/ALU/_340_ ) );
NAND2_X1 \EXU/ALU/_650_ ( .A1(\EXU/ALU/_144_ ), .A2(\EXU/ALU/_112_ ), .ZN(\EXU/ALU/_341_ ) );
NAND4_X1 \EXU/ALU/_651_ ( .A1(\EXU/ALU/_340_ ), .A2(fanout_net_15 ), .A3(\EXU/ALU/_332_ ), .A4(\EXU/ALU/_341_ ), .ZN(\EXU/ALU/_342_ ) );
NAND4_X1 \EXU/ALU/_652_ ( .A1(\EXU/ALU/_264_ ), .A2(fanout_net_12 ), .A3(fanout_net_13 ), .A4(\EXU/ALU/_144_ ), .ZN(\EXU/ALU/_343_ ) );
AND2_X1 \EXU/ALU/_653_ ( .A1(\EXU/ALU/_342_ ), .A2(\EXU/ALU/_343_ ), .ZN(\EXU/ALU/_344_ ) );
NAND3_X1 \EXU/ALU/_654_ ( .A1(\EXU/ALU/_285_ ), .A2(\EXU/ALU/_286_ ), .A3(\EXU/ALU/_011_ ), .ZN(\EXU/ALU/_345_ ) );
AOI22_X1 \EXU/ALU/_655_ ( .A1(\EXU/ALU/_276_ ), .A2(\EXU/ALU/_340_ ), .B1(\EXU/ALU/_048_ ), .B2(\EXU/ALU/_277_ ), .ZN(\EXU/ALU/_346_ ) );
NAND4_X1 \EXU/ALU/_656_ ( .A1(\EXU/ALU/_289_ ), .A2(fanout_net_15 ), .A3(\EXU/ALU/_144_ ), .A4(\EXU/ALU/_112_ ), .ZN(\EXU/ALU/_347_ ) );
NAND4_X1 \EXU/ALU/_657_ ( .A1(\EXU/ALU/_344_ ), .A2(\EXU/ALU/_345_ ), .A3(\EXU/ALU/_346_ ), .A4(\EXU/ALU/_347_ ), .ZN(\EXU/ALU/_080_ ) );
OR2_X1 \EXU/ALU/_658_ ( .A1(\EXU/ALU/_145_ ), .A2(\EXU/ALU/_113_ ), .ZN(\EXU/ALU/_348_ ) );
NAND2_X1 \EXU/ALU/_659_ ( .A1(\EXU/ALU/_145_ ), .A2(\EXU/ALU/_113_ ), .ZN(\EXU/ALU/_349_ ) );
NAND4_X1 \EXU/ALU/_660_ ( .A1(\EXU/ALU/_348_ ), .A2(fanout_net_15 ), .A3(\EXU/ALU/_332_ ), .A4(\EXU/ALU/_349_ ), .ZN(\EXU/ALU/_350_ ) );
BUF_X8 \EXU/ALU/_661_ ( .A(\EXU/ALU/_174_ ), .Z(\EXU/ALU/_351_ ) );
NAND4_X1 \EXU/ALU/_662_ ( .A1(\EXU/ALU/_351_ ), .A2(fanout_net_12 ), .A3(fanout_net_13 ), .A4(\EXU/ALU/_145_ ), .ZN(\EXU/ALU/_352_ ) );
AND2_X1 \EXU/ALU/_663_ ( .A1(\EXU/ALU/_350_ ), .A2(\EXU/ALU/_352_ ), .ZN(\EXU/ALU/_353_ ) );
NAND3_X1 \EXU/ALU/_664_ ( .A1(\EXU/ALU/_285_ ), .A2(\EXU/ALU/_286_ ), .A3(\EXU/ALU/_012_ ), .ZN(\EXU/ALU/_354_ ) );
AOI22_X1 \EXU/ALU/_665_ ( .A1(\EXU/ALU/_276_ ), .A2(\EXU/ALU/_348_ ), .B1(\EXU/ALU/_049_ ), .B2(\EXU/ALU/_277_ ), .ZN(\EXU/ALU/_355_ ) );
NAND4_X1 \EXU/ALU/_666_ ( .A1(\EXU/ALU/_289_ ), .A2(fanout_net_15 ), .A3(\EXU/ALU/_145_ ), .A4(\EXU/ALU/_113_ ), .ZN(\EXU/ALU/_356_ ) );
NAND4_X1 \EXU/ALU/_667_ ( .A1(\EXU/ALU/_353_ ), .A2(\EXU/ALU/_354_ ), .A3(\EXU/ALU/_355_ ), .A4(\EXU/ALU/_356_ ), .ZN(\EXU/ALU/_081_ ) );
OR2_X1 \EXU/ALU/_668_ ( .A1(\EXU/ALU/_147_ ), .A2(\EXU/ALU/_115_ ), .ZN(\EXU/ALU/_357_ ) );
NAND2_X1 \EXU/ALU/_669_ ( .A1(\EXU/ALU/_147_ ), .A2(\EXU/ALU/_115_ ), .ZN(\EXU/ALU/_358_ ) );
NAND4_X1 \EXU/ALU/_670_ ( .A1(\EXU/ALU/_357_ ), .A2(fanout_net_15 ), .A3(\EXU/ALU/_332_ ), .A4(\EXU/ALU/_358_ ), .ZN(\EXU/ALU/_359_ ) );
NAND4_X1 \EXU/ALU/_671_ ( .A1(\EXU/ALU/_351_ ), .A2(fanout_net_12 ), .A3(fanout_net_13 ), .A4(\EXU/ALU/_147_ ), .ZN(\EXU/ALU/_360_ ) );
AND2_X1 \EXU/ALU/_672_ ( .A1(\EXU/ALU/_359_ ), .A2(\EXU/ALU/_360_ ), .ZN(\EXU/ALU/_361_ ) );
NAND3_X1 \EXU/ALU/_673_ ( .A1(\EXU/ALU/_285_ ), .A2(\EXU/ALU/_286_ ), .A3(\EXU/ALU/_014_ ), .ZN(\EXU/ALU/_362_ ) );
BUF_X4 \EXU/ALU/_674_ ( .A(\EXU/ALU/_182_ ), .Z(\EXU/ALU/_363_ ) );
BUF_X4 \EXU/ALU/_675_ ( .A(\EXU/ALU/_189_ ), .Z(\EXU/ALU/_364_ ) );
AOI22_X1 \EXU/ALU/_676_ ( .A1(\EXU/ALU/_363_ ), .A2(\EXU/ALU/_357_ ), .B1(\EXU/ALU/_051_ ), .B2(\EXU/ALU/_364_ ), .ZN(\EXU/ALU/_365_ ) );
NAND4_X1 \EXU/ALU/_677_ ( .A1(\EXU/ALU/_289_ ), .A2(fanout_net_15 ), .A3(\EXU/ALU/_147_ ), .A4(\EXU/ALU/_115_ ), .ZN(\EXU/ALU/_366_ ) );
NAND4_X1 \EXU/ALU/_678_ ( .A1(\EXU/ALU/_361_ ), .A2(\EXU/ALU/_362_ ), .A3(\EXU/ALU/_365_ ), .A4(\EXU/ALU/_366_ ), .ZN(\EXU/ALU/_083_ ) );
OR2_X1 \EXU/ALU/_679_ ( .A1(\EXU/ALU/_148_ ), .A2(\EXU/ALU/_116_ ), .ZN(\EXU/ALU/_367_ ) );
NAND2_X1 \EXU/ALU/_680_ ( .A1(\EXU/ALU/_148_ ), .A2(\EXU/ALU/_116_ ), .ZN(\EXU/ALU/_368_ ) );
NAND4_X1 \EXU/ALU/_681_ ( .A1(\EXU/ALU/_367_ ), .A2(fanout_net_15 ), .A3(\EXU/ALU/_332_ ), .A4(\EXU/ALU/_368_ ), .ZN(\EXU/ALU/_369_ ) );
NAND4_X1 \EXU/ALU/_682_ ( .A1(\EXU/ALU/_351_ ), .A2(fanout_net_12 ), .A3(fanout_net_13 ), .A4(\EXU/ALU/_148_ ), .ZN(\EXU/ALU/_370_ ) );
AND2_X1 \EXU/ALU/_683_ ( .A1(\EXU/ALU/_369_ ), .A2(\EXU/ALU/_370_ ), .ZN(\EXU/ALU/_371_ ) );
BUF_X4 \EXU/ALU/_684_ ( .A(\EXU/ALU/_193_ ), .Z(\EXU/ALU/_372_ ) );
BUF_X4 \EXU/ALU/_685_ ( .A(\EXU/ALU/_174_ ), .Z(\EXU/ALU/_373_ ) );
NAND3_X1 \EXU/ALU/_686_ ( .A1(\EXU/ALU/_372_ ), .A2(\EXU/ALU/_373_ ), .A3(\EXU/ALU/_015_ ), .ZN(\EXU/ALU/_374_ ) );
AOI22_X1 \EXU/ALU/_687_ ( .A1(\EXU/ALU/_363_ ), .A2(\EXU/ALU/_367_ ), .B1(\EXU/ALU/_052_ ), .B2(\EXU/ALU/_364_ ), .ZN(\EXU/ALU/_375_ ) );
BUF_X4 \EXU/ALU/_688_ ( .A(\EXU/ALU/_185_ ), .Z(\EXU/ALU/_376_ ) );
NAND4_X1 \EXU/ALU/_689_ ( .A1(\EXU/ALU/_376_ ), .A2(fanout_net_15 ), .A3(\EXU/ALU/_148_ ), .A4(\EXU/ALU/_116_ ), .ZN(\EXU/ALU/_377_ ) );
NAND4_X1 \EXU/ALU/_690_ ( .A1(\EXU/ALU/_371_ ), .A2(\EXU/ALU/_374_ ), .A3(\EXU/ALU/_375_ ), .A4(\EXU/ALU/_377_ ), .ZN(\EXU/ALU/_084_ ) );
OR2_X1 \EXU/ALU/_691_ ( .A1(\EXU/ALU/_149_ ), .A2(\EXU/ALU/_117_ ), .ZN(\EXU/ALU/_378_ ) );
NAND2_X1 \EXU/ALU/_692_ ( .A1(\EXU/ALU/_149_ ), .A2(\EXU/ALU/_117_ ), .ZN(\EXU/ALU/_379_ ) );
NAND4_X1 \EXU/ALU/_693_ ( .A1(\EXU/ALU/_378_ ), .A2(fanout_net_15 ), .A3(\EXU/ALU/_332_ ), .A4(\EXU/ALU/_379_ ), .ZN(\EXU/ALU/_380_ ) );
NAND4_X1 \EXU/ALU/_694_ ( .A1(\EXU/ALU/_351_ ), .A2(fanout_net_12 ), .A3(fanout_net_13 ), .A4(\EXU/ALU/_149_ ), .ZN(\EXU/ALU/_381_ ) );
AND2_X1 \EXU/ALU/_695_ ( .A1(\EXU/ALU/_380_ ), .A2(\EXU/ALU/_381_ ), .ZN(\EXU/ALU/_382_ ) );
NAND3_X1 \EXU/ALU/_696_ ( .A1(\EXU/ALU/_372_ ), .A2(\EXU/ALU/_373_ ), .A3(\EXU/ALU/_016_ ), .ZN(\EXU/ALU/_383_ ) );
AOI22_X1 \EXU/ALU/_697_ ( .A1(\EXU/ALU/_363_ ), .A2(\EXU/ALU/_378_ ), .B1(\EXU/ALU/_053_ ), .B2(\EXU/ALU/_364_ ), .ZN(\EXU/ALU/_384_ ) );
NAND4_X1 \EXU/ALU/_698_ ( .A1(\EXU/ALU/_376_ ), .A2(fanout_net_15 ), .A3(\EXU/ALU/_149_ ), .A4(\EXU/ALU/_117_ ), .ZN(\EXU/ALU/_385_ ) );
NAND4_X1 \EXU/ALU/_699_ ( .A1(\EXU/ALU/_382_ ), .A2(\EXU/ALU/_383_ ), .A3(\EXU/ALU/_384_ ), .A4(\EXU/ALU/_385_ ), .ZN(\EXU/ALU/_085_ ) );
OR2_X1 \EXU/ALU/_700_ ( .A1(\EXU/ALU/_150_ ), .A2(\EXU/ALU/_118_ ), .ZN(\EXU/ALU/_386_ ) );
NAND2_X1 \EXU/ALU/_701_ ( .A1(\EXU/ALU/_150_ ), .A2(\EXU/ALU/_118_ ), .ZN(\EXU/ALU/_387_ ) );
NAND4_X1 \EXU/ALU/_702_ ( .A1(\EXU/ALU/_386_ ), .A2(fanout_net_15 ), .A3(\EXU/ALU/_332_ ), .A4(\EXU/ALU/_387_ ), .ZN(\EXU/ALU/_388_ ) );
NAND4_X1 \EXU/ALU/_703_ ( .A1(\EXU/ALU/_351_ ), .A2(fanout_net_12 ), .A3(fanout_net_13 ), .A4(\EXU/ALU/_150_ ), .ZN(\EXU/ALU/_389_ ) );
AND2_X1 \EXU/ALU/_704_ ( .A1(\EXU/ALU/_388_ ), .A2(\EXU/ALU/_389_ ), .ZN(\EXU/ALU/_390_ ) );
NAND3_X1 \EXU/ALU/_705_ ( .A1(\EXU/ALU/_372_ ), .A2(\EXU/ALU/_373_ ), .A3(\EXU/ALU/_017_ ), .ZN(\EXU/ALU/_391_ ) );
AOI22_X1 \EXU/ALU/_706_ ( .A1(\EXU/ALU/_363_ ), .A2(\EXU/ALU/_386_ ), .B1(\EXU/ALU/_054_ ), .B2(\EXU/ALU/_364_ ), .ZN(\EXU/ALU/_392_ ) );
NAND4_X1 \EXU/ALU/_707_ ( .A1(\EXU/ALU/_376_ ), .A2(fanout_net_15 ), .A3(\EXU/ALU/_150_ ), .A4(\EXU/ALU/_118_ ), .ZN(\EXU/ALU/_393_ ) );
NAND4_X1 \EXU/ALU/_708_ ( .A1(\EXU/ALU/_390_ ), .A2(\EXU/ALU/_391_ ), .A3(\EXU/ALU/_392_ ), .A4(\EXU/ALU/_393_ ), .ZN(\EXU/ALU/_086_ ) );
OR2_X1 \EXU/ALU/_709_ ( .A1(\EXU/ALU/_151_ ), .A2(\EXU/ALU/_119_ ), .ZN(\EXU/ALU/_394_ ) );
NAND2_X1 \EXU/ALU/_710_ ( .A1(\EXU/ALU/_151_ ), .A2(\EXU/ALU/_119_ ), .ZN(\EXU/ALU/_395_ ) );
NAND4_X1 \EXU/ALU/_711_ ( .A1(\EXU/ALU/_394_ ), .A2(fanout_net_15 ), .A3(\EXU/ALU/_332_ ), .A4(\EXU/ALU/_395_ ), .ZN(\EXU/ALU/_396_ ) );
NAND4_X1 \EXU/ALU/_712_ ( .A1(\EXU/ALU/_351_ ), .A2(fanout_net_12 ), .A3(fanout_net_13 ), .A4(\EXU/ALU/_151_ ), .ZN(\EXU/ALU/_397_ ) );
AND2_X2 \EXU/ALU/_713_ ( .A1(\EXU/ALU/_396_ ), .A2(\EXU/ALU/_397_ ), .ZN(\EXU/ALU/_398_ ) );
NAND3_X1 \EXU/ALU/_714_ ( .A1(\EXU/ALU/_372_ ), .A2(\EXU/ALU/_373_ ), .A3(\EXU/ALU/_018_ ), .ZN(\EXU/ALU/_399_ ) );
AOI22_X1 \EXU/ALU/_715_ ( .A1(\EXU/ALU/_363_ ), .A2(\EXU/ALU/_394_ ), .B1(\EXU/ALU/_055_ ), .B2(\EXU/ALU/_364_ ), .ZN(\EXU/ALU/_400_ ) );
NAND4_X1 \EXU/ALU/_716_ ( .A1(\EXU/ALU/_376_ ), .A2(fanout_net_15 ), .A3(\EXU/ALU/_151_ ), .A4(\EXU/ALU/_119_ ), .ZN(\EXU/ALU/_401_ ) );
NAND4_X1 \EXU/ALU/_717_ ( .A1(\EXU/ALU/_398_ ), .A2(\EXU/ALU/_399_ ), .A3(\EXU/ALU/_400_ ), .A4(\EXU/ALU/_401_ ), .ZN(\EXU/ALU/_087_ ) );
OR2_X1 \EXU/ALU/_718_ ( .A1(\EXU/ALU/_152_ ), .A2(\EXU/ALU/_120_ ), .ZN(\EXU/ALU/_402_ ) );
NAND2_X1 \EXU/ALU/_719_ ( .A1(\EXU/ALU/_152_ ), .A2(\EXU/ALU/_120_ ), .ZN(\EXU/ALU/_403_ ) );
NAND4_X1 \EXU/ALU/_720_ ( .A1(\EXU/ALU/_402_ ), .A2(fanout_net_15 ), .A3(\EXU/ALU/_332_ ), .A4(\EXU/ALU/_403_ ), .ZN(\EXU/ALU/_404_ ) );
NAND4_X1 \EXU/ALU/_721_ ( .A1(\EXU/ALU/_351_ ), .A2(fanout_net_12 ), .A3(fanout_net_13 ), .A4(\EXU/ALU/_152_ ), .ZN(\EXU/ALU/_405_ ) );
AND2_X2 \EXU/ALU/_722_ ( .A1(\EXU/ALU/_404_ ), .A2(\EXU/ALU/_405_ ), .ZN(\EXU/ALU/_406_ ) );
NAND3_X1 \EXU/ALU/_723_ ( .A1(\EXU/ALU/_372_ ), .A2(\EXU/ALU/_373_ ), .A3(\EXU/ALU/_019_ ), .ZN(\EXU/ALU/_407_ ) );
AOI22_X1 \EXU/ALU/_724_ ( .A1(\EXU/ALU/_363_ ), .A2(\EXU/ALU/_402_ ), .B1(\EXU/ALU/_056_ ), .B2(\EXU/ALU/_364_ ), .ZN(\EXU/ALU/_408_ ) );
NAND4_X1 \EXU/ALU/_725_ ( .A1(\EXU/ALU/_376_ ), .A2(fanout_net_15 ), .A3(\EXU/ALU/_152_ ), .A4(\EXU/ALU/_120_ ), .ZN(\EXU/ALU/_409_ ) );
NAND4_X1 \EXU/ALU/_726_ ( .A1(\EXU/ALU/_406_ ), .A2(\EXU/ALU/_407_ ), .A3(\EXU/ALU/_408_ ), .A4(\EXU/ALU/_409_ ), .ZN(\EXU/ALU/_088_ ) );
OR2_X1 \EXU/ALU/_727_ ( .A1(\EXU/ALU/_153_ ), .A2(\EXU/ALU/_121_ ), .ZN(\EXU/ALU/_410_ ) );
NAND2_X1 \EXU/ALU/_728_ ( .A1(\EXU/ALU/_153_ ), .A2(\EXU/ALU/_121_ ), .ZN(\EXU/ALU/_411_ ) );
NAND4_X1 \EXU/ALU/_729_ ( .A1(\EXU/ALU/_410_ ), .A2(fanout_net_15 ), .A3(\EXU/ALU/_332_ ), .A4(\EXU/ALU/_411_ ), .ZN(\EXU/ALU/_412_ ) );
NAND4_X1 \EXU/ALU/_730_ ( .A1(\EXU/ALU/_351_ ), .A2(fanout_net_12 ), .A3(\EXU/ALU/_035_ ), .A4(\EXU/ALU/_153_ ), .ZN(\EXU/ALU/_413_ ) );
AND2_X2 \EXU/ALU/_731_ ( .A1(\EXU/ALU/_412_ ), .A2(\EXU/ALU/_413_ ), .ZN(\EXU/ALU/_414_ ) );
NAND3_X1 \EXU/ALU/_732_ ( .A1(\EXU/ALU/_372_ ), .A2(\EXU/ALU/_373_ ), .A3(\EXU/ALU/_020_ ), .ZN(\EXU/ALU/_415_ ) );
AOI22_X1 \EXU/ALU/_733_ ( .A1(\EXU/ALU/_363_ ), .A2(\EXU/ALU/_410_ ), .B1(\EXU/ALU/_057_ ), .B2(\EXU/ALU/_364_ ), .ZN(\EXU/ALU/_416_ ) );
NAND4_X1 \EXU/ALU/_734_ ( .A1(\EXU/ALU/_376_ ), .A2(fanout_net_15 ), .A3(\EXU/ALU/_153_ ), .A4(\EXU/ALU/_121_ ), .ZN(\EXU/ALU/_417_ ) );
NAND4_X1 \EXU/ALU/_735_ ( .A1(\EXU/ALU/_414_ ), .A2(\EXU/ALU/_415_ ), .A3(\EXU/ALU/_416_ ), .A4(\EXU/ALU/_417_ ), .ZN(\EXU/ALU/_089_ ) );
OR2_X1 \EXU/ALU/_736_ ( .A1(\EXU/ALU/_154_ ), .A2(\EXU/ALU/_122_ ), .ZN(\EXU/ALU/_418_ ) );
NAND2_X1 \EXU/ALU/_737_ ( .A1(\EXU/ALU/_154_ ), .A2(\EXU/ALU/_122_ ), .ZN(\EXU/ALU/_419_ ) );
NAND4_X1 \EXU/ALU/_738_ ( .A1(\EXU/ALU/_418_ ), .A2(fanout_net_15 ), .A3(\EXU/ALU/_178_ ), .A4(\EXU/ALU/_419_ ), .ZN(\EXU/ALU/_420_ ) );
NAND4_X1 \EXU/ALU/_739_ ( .A1(\EXU/ALU/_351_ ), .A2(fanout_net_12 ), .A3(\EXU/ALU/_035_ ), .A4(\EXU/ALU/_154_ ), .ZN(\EXU/ALU/_421_ ) );
AND2_X1 \EXU/ALU/_740_ ( .A1(\EXU/ALU/_420_ ), .A2(\EXU/ALU/_421_ ), .ZN(\EXU/ALU/_422_ ) );
NAND3_X1 \EXU/ALU/_741_ ( .A1(\EXU/ALU/_372_ ), .A2(\EXU/ALU/_373_ ), .A3(\EXU/ALU/_021_ ), .ZN(\EXU/ALU/_423_ ) );
AOI22_X1 \EXU/ALU/_742_ ( .A1(\EXU/ALU/_363_ ), .A2(\EXU/ALU/_418_ ), .B1(\EXU/ALU/_058_ ), .B2(\EXU/ALU/_364_ ), .ZN(\EXU/ALU/_424_ ) );
NAND4_X1 \EXU/ALU/_743_ ( .A1(\EXU/ALU/_376_ ), .A2(fanout_net_15 ), .A3(\EXU/ALU/_154_ ), .A4(\EXU/ALU/_122_ ), .ZN(\EXU/ALU/_425_ ) );
NAND4_X1 \EXU/ALU/_744_ ( .A1(\EXU/ALU/_422_ ), .A2(\EXU/ALU/_423_ ), .A3(\EXU/ALU/_424_ ), .A4(\EXU/ALU/_425_ ), .ZN(\EXU/ALU/_090_ ) );
OR2_X1 \EXU/ALU/_745_ ( .A1(\EXU/ALU/_155_ ), .A2(\EXU/ALU/_123_ ), .ZN(\EXU/ALU/_426_ ) );
NAND2_X1 \EXU/ALU/_746_ ( .A1(\EXU/ALU/_155_ ), .A2(\EXU/ALU/_123_ ), .ZN(\EXU/ALU/_427_ ) );
NAND4_X1 \EXU/ALU/_747_ ( .A1(\EXU/ALU/_426_ ), .A2(fanout_net_15 ), .A3(\EXU/ALU/_178_ ), .A4(\EXU/ALU/_427_ ), .ZN(\EXU/ALU/_428_ ) );
NAND4_X1 \EXU/ALU/_748_ ( .A1(\EXU/ALU/_351_ ), .A2(\EXU/ALU/_034_ ), .A3(\EXU/ALU/_035_ ), .A4(\EXU/ALU/_155_ ), .ZN(\EXU/ALU/_429_ ) );
AND2_X1 \EXU/ALU/_749_ ( .A1(\EXU/ALU/_428_ ), .A2(\EXU/ALU/_429_ ), .ZN(\EXU/ALU/_430_ ) );
NAND3_X1 \EXU/ALU/_750_ ( .A1(\EXU/ALU/_372_ ), .A2(\EXU/ALU/_373_ ), .A3(\EXU/ALU/_022_ ), .ZN(\EXU/ALU/_431_ ) );
AOI22_X1 \EXU/ALU/_751_ ( .A1(\EXU/ALU/_363_ ), .A2(\EXU/ALU/_426_ ), .B1(\EXU/ALU/_059_ ), .B2(\EXU/ALU/_364_ ), .ZN(\EXU/ALU/_432_ ) );
NAND4_X1 \EXU/ALU/_752_ ( .A1(\EXU/ALU/_376_ ), .A2(fanout_net_15 ), .A3(\EXU/ALU/_155_ ), .A4(\EXU/ALU/_123_ ), .ZN(\EXU/ALU/_433_ ) );
NAND4_X1 \EXU/ALU/_753_ ( .A1(\EXU/ALU/_430_ ), .A2(\EXU/ALU/_431_ ), .A3(\EXU/ALU/_432_ ), .A4(\EXU/ALU/_433_ ), .ZN(\EXU/ALU/_091_ ) );
OR2_X1 \EXU/ALU/_754_ ( .A1(\EXU/ALU/_156_ ), .A2(\EXU/ALU/_124_ ), .ZN(\EXU/ALU/_434_ ) );
NAND2_X1 \EXU/ALU/_755_ ( .A1(\EXU/ALU/_156_ ), .A2(\EXU/ALU/_124_ ), .ZN(\EXU/ALU/_435_ ) );
NAND4_X1 \EXU/ALU/_756_ ( .A1(\EXU/ALU/_434_ ), .A2(fanout_net_15 ), .A3(\EXU/ALU/_178_ ), .A4(\EXU/ALU/_435_ ), .ZN(\EXU/ALU/_436_ ) );
NAND4_X1 \EXU/ALU/_757_ ( .A1(\EXU/ALU/_174_ ), .A2(\EXU/ALU/_034_ ), .A3(\EXU/ALU/_035_ ), .A4(\EXU/ALU/_156_ ), .ZN(\EXU/ALU/_437_ ) );
AND2_X1 \EXU/ALU/_758_ ( .A1(\EXU/ALU/_436_ ), .A2(\EXU/ALU/_437_ ), .ZN(\EXU/ALU/_438_ ) );
NAND3_X1 \EXU/ALU/_759_ ( .A1(\EXU/ALU/_372_ ), .A2(\EXU/ALU/_373_ ), .A3(\EXU/ALU/_023_ ), .ZN(\EXU/ALU/_439_ ) );
AOI22_X1 \EXU/ALU/_760_ ( .A1(\EXU/ALU/_363_ ), .A2(\EXU/ALU/_434_ ), .B1(\EXU/ALU/_060_ ), .B2(\EXU/ALU/_364_ ), .ZN(\EXU/ALU/_440_ ) );
NAND4_X1 \EXU/ALU/_761_ ( .A1(\EXU/ALU/_376_ ), .A2(fanout_net_15 ), .A3(\EXU/ALU/_156_ ), .A4(\EXU/ALU/_124_ ), .ZN(\EXU/ALU/_441_ ) );
NAND4_X1 \EXU/ALU/_762_ ( .A1(\EXU/ALU/_438_ ), .A2(\EXU/ALU/_439_ ), .A3(\EXU/ALU/_440_ ), .A4(\EXU/ALU/_441_ ), .ZN(\EXU/ALU/_092_ ) );
OR2_X1 \EXU/ALU/_763_ ( .A1(\EXU/ALU/_158_ ), .A2(\EXU/ALU/_126_ ), .ZN(\EXU/ALU/_442_ ) );
NAND2_X1 \EXU/ALU/_764_ ( .A1(\EXU/ALU/_158_ ), .A2(\EXU/ALU/_126_ ), .ZN(\EXU/ALU/_443_ ) );
NAND4_X1 \EXU/ALU/_765_ ( .A1(\EXU/ALU/_442_ ), .A2(\EXU/ALU/_036_ ), .A3(\EXU/ALU/_178_ ), .A4(\EXU/ALU/_443_ ), .ZN(\EXU/ALU/_444_ ) );
NAND4_X1 \EXU/ALU/_766_ ( .A1(\EXU/ALU/_174_ ), .A2(\EXU/ALU/_034_ ), .A3(\EXU/ALU/_035_ ), .A4(\EXU/ALU/_158_ ), .ZN(\EXU/ALU/_445_ ) );
AND2_X1 \EXU/ALU/_767_ ( .A1(\EXU/ALU/_444_ ), .A2(\EXU/ALU/_445_ ), .ZN(\EXU/ALU/_446_ ) );
NAND3_X1 \EXU/ALU/_768_ ( .A1(\EXU/ALU/_372_ ), .A2(\EXU/ALU/_373_ ), .A3(\EXU/ALU/_025_ ), .ZN(\EXU/ALU/_447_ ) );
AOI22_X1 \EXU/ALU/_769_ ( .A1(\EXU/ALU/_182_ ), .A2(\EXU/ALU/_442_ ), .B1(\EXU/ALU/_062_ ), .B2(\EXU/ALU/_189_ ), .ZN(\EXU/ALU/_448_ ) );
NAND4_X1 \EXU/ALU/_770_ ( .A1(\EXU/ALU/_376_ ), .A2(\EXU/ALU/_036_ ), .A3(\EXU/ALU/_158_ ), .A4(\EXU/ALU/_126_ ), .ZN(\EXU/ALU/_449_ ) );
NAND4_X1 \EXU/ALU/_771_ ( .A1(\EXU/ALU/_446_ ), .A2(\EXU/ALU/_447_ ), .A3(\EXU/ALU/_448_ ), .A4(\EXU/ALU/_449_ ), .ZN(\EXU/ALU/_094_ ) );
OR2_X1 \EXU/ALU/_772_ ( .A1(\EXU/ALU/_159_ ), .A2(\EXU/ALU/_127_ ), .ZN(\EXU/ALU/_450_ ) );
NAND2_X1 \EXU/ALU/_773_ ( .A1(\EXU/ALU/_159_ ), .A2(\EXU/ALU/_127_ ), .ZN(\EXU/ALU/_451_ ) );
NAND4_X1 \EXU/ALU/_774_ ( .A1(\EXU/ALU/_450_ ), .A2(\EXU/ALU/_036_ ), .A3(\EXU/ALU/_178_ ), .A4(\EXU/ALU/_451_ ), .ZN(\EXU/ALU/_452_ ) );
NAND4_X1 \EXU/ALU/_775_ ( .A1(\EXU/ALU/_174_ ), .A2(\EXU/ALU/_034_ ), .A3(\EXU/ALU/_035_ ), .A4(\EXU/ALU/_159_ ), .ZN(\EXU/ALU/_453_ ) );
AND2_X1 \EXU/ALU/_776_ ( .A1(\EXU/ALU/_452_ ), .A2(\EXU/ALU/_453_ ), .ZN(\EXU/ALU/_454_ ) );
NAND3_X1 \EXU/ALU/_777_ ( .A1(\EXU/ALU/_193_ ), .A2(\EXU/ALU/_026_ ), .A3(\EXU/ALU/_186_ ), .ZN(\EXU/ALU/_455_ ) );
AOI22_X1 \EXU/ALU/_778_ ( .A1(\EXU/ALU/_182_ ), .A2(\EXU/ALU/_450_ ), .B1(\EXU/ALU/_063_ ), .B2(\EXU/ALU/_189_ ), .ZN(\EXU/ALU/_456_ ) );
NAND4_X1 \EXU/ALU/_779_ ( .A1(\EXU/ALU/_185_ ), .A2(\EXU/ALU/_036_ ), .A3(\EXU/ALU/_159_ ), .A4(\EXU/ALU/_127_ ), .ZN(\EXU/ALU/_457_ ) );
NAND4_X1 \EXU/ALU/_780_ ( .A1(\EXU/ALU/_454_ ), .A2(\EXU/ALU/_455_ ), .A3(\EXU/ALU/_456_ ), .A4(\EXU/ALU/_457_ ), .ZN(\EXU/ALU/_095_ ) );
BUF_X1 \EXU/ALU/_781_ ( .A(\EXU/ALU/_adder_io_result [31] ), .Z(\EXU/ALU/_026_ ) );
BUF_X1 \EXU/ALU/_782_ ( .A(\EXU/ALU/_adder_io_overflow ), .Z(\EXU/ALU/_001_ ) );
BUF_X1 \EXU/ALU/_783_ ( .A(\EXU/ALU/_aluControl_io_isSub ), .Z(\EXU/ALU/_037_ ) );
BUF_X1 \EXU/ALU/_784_ ( .A(\EXU/ALU/_adder_io_carry ), .Z(\EXU/ALU/_000_ ) );
BUF_X1 \EXU/ALU/_785_ ( .A(\EXU/ALU/_aluControl_io_isUnsigned ), .Z(\EXU/ALU/_038_ ) );
BUF_X1 \EXU/ALU/_786_ ( .A(\EXU/ALU/_167_ ), .Z(\EXU/_ALU_io_less ) );
BUF_X1 \EXU/ALU/_787_ ( .A(\EXU/casez_tmp_0 [0] ), .Z(\EXU/ALU/_135_ ) );
BUF_X1 \EXU/ALU/_788_ ( .A(\EXU/_0000_ ), .Z(\EXU/ALU/_103_ ) );
BUF_X1 \EXU/ALU/_789_ ( .A(\EXU/ALU/_aluControl_io_aluSel [0] ), .Z(\EXU/ALU/_034_ ) );
BUF_X1 \EXU/ALU/_790_ ( .A(\EXU/ALU/_aluControl_io_aluSel [1] ), .Z(\EXU/ALU/_035_ ) );
BUF_X1 \EXU/ALU/_791_ ( .A(\EXU/ALU/_aluControl_io_aluSel [2] ), .Z(\EXU/ALU/_036_ ) );
BUF_X1 \EXU/ALU/_792_ ( .A(\EXU/ALU/_barrelShift_io_out [0] ), .Z(\EXU/ALU/_039_ ) );
BUF_X1 \EXU/ALU/_793_ ( .A(\EXU/ALU/_adder_io_result [0] ), .Z(\EXU/ALU/_002_ ) );
BUF_X1 \EXU/ALU/_794_ ( .A(\EXU/ALU/_071_ ), .Z(\_EXU_io_LSUIn_bits_raddr [0] ) );
BUF_X1 \EXU/ALU/_795_ ( .A(\EXU/casez_tmp_0 [1] ), .Z(\EXU/ALU/_146_ ) );
BUF_X1 \EXU/ALU/_796_ ( .A(\EXU/_0011_ ), .Z(\EXU/ALU/_114_ ) );
BUF_X1 \EXU/ALU/_797_ ( .A(\EXU/ALU/_barrelShift_io_out [1] ), .Z(\EXU/ALU/_050_ ) );
BUF_X1 \EXU/ALU/_798_ ( .A(\EXU/ALU/_adder_io_result [1] ), .Z(\EXU/ALU/_013_ ) );
BUF_X1 \EXU/ALU/_799_ ( .A(\EXU/ALU/_082_ ), .Z(\_EXU_io_LSUIn_bits_raddr [1] ) );
BUF_X1 \EXU/ALU/_800_ ( .A(\EXU/casez_tmp_0 [2] ), .Z(\EXU/ALU/_157_ ) );
BUF_X1 \EXU/ALU/_801_ ( .A(\EXU/_0022_ ), .Z(\EXU/ALU/_125_ ) );
BUF_X1 \EXU/ALU/_802_ ( .A(\EXU/ALU/_barrelShift_io_out [2] ), .Z(\EXU/ALU/_061_ ) );
BUF_X1 \EXU/ALU/_803_ ( .A(\EXU/ALU/_adder_io_result [2] ), .Z(\EXU/ALU/_024_ ) );
BUF_X1 \EXU/ALU/_804_ ( .A(\EXU/ALU/_093_ ), .Z(\_EXU_io_LSUIn_bits_raddr [2] ) );
BUF_X1 \EXU/ALU/_805_ ( .A(\EXU/casez_tmp_0 [3] ), .Z(\EXU/ALU/_160_ ) );
BUF_X1 \EXU/ALU/_806_ ( .A(\EXU/_0025_ ), .Z(\EXU/ALU/_128_ ) );
BUF_X1 \EXU/ALU/_807_ ( .A(\EXU/ALU/_barrelShift_io_out [3] ), .Z(\EXU/ALU/_064_ ) );
BUF_X1 \EXU/ALU/_808_ ( .A(\EXU/ALU/_adder_io_result [3] ), .Z(\EXU/ALU/_027_ ) );
BUF_X1 \EXU/ALU/_809_ ( .A(\EXU/ALU/_096_ ), .Z(\_EXU_io_LSUIn_bits_raddr [3] ) );
BUF_X1 \EXU/ALU/_810_ ( .A(\EXU/casez_tmp_0 [4] ), .Z(\EXU/ALU/_161_ ) );
BUF_X1 \EXU/ALU/_811_ ( .A(\EXU/_0026_ ), .Z(\EXU/ALU/_129_ ) );
BUF_X1 \EXU/ALU/_812_ ( .A(\EXU/ALU/_barrelShift_io_out [4] ), .Z(\EXU/ALU/_065_ ) );
BUF_X1 \EXU/ALU/_813_ ( .A(\EXU/ALU/_adder_io_result [4] ), .Z(\EXU/ALU/_028_ ) );
BUF_X1 \EXU/ALU/_814_ ( .A(\EXU/ALU/_097_ ), .Z(\_EXU_io_LSUIn_bits_raddr [4] ) );
BUF_X1 \EXU/ALU/_815_ ( .A(\EXU/casez_tmp_0 [5] ), .Z(\EXU/ALU/_162_ ) );
BUF_X1 \EXU/ALU/_816_ ( .A(\EXU/_0027_ ), .Z(\EXU/ALU/_130_ ) );
BUF_X1 \EXU/ALU/_817_ ( .A(\EXU/ALU/_barrelShift_io_out [5] ), .Z(\EXU/ALU/_066_ ) );
BUF_X1 \EXU/ALU/_818_ ( .A(\EXU/ALU/_adder_io_result [5] ), .Z(\EXU/ALU/_029_ ) );
BUF_X1 \EXU/ALU/_819_ ( .A(\EXU/ALU/_098_ ), .Z(\_EXU_io_LSUIn_bits_raddr [5] ) );
BUF_X1 \EXU/ALU/_820_ ( .A(\EXU/casez_tmp_0 [6] ), .Z(\EXU/ALU/_163_ ) );
BUF_X1 \EXU/ALU/_821_ ( .A(\EXU/_0028_ ), .Z(\EXU/ALU/_131_ ) );
BUF_X1 \EXU/ALU/_822_ ( .A(\EXU/ALU/_barrelShift_io_out [6] ), .Z(\EXU/ALU/_067_ ) );
BUF_X1 \EXU/ALU/_823_ ( .A(\EXU/ALU/_adder_io_result [6] ), .Z(\EXU/ALU/_030_ ) );
BUF_X1 \EXU/ALU/_824_ ( .A(\EXU/ALU/_099_ ), .Z(\_EXU_io_LSUIn_bits_raddr [6] ) );
BUF_X1 \EXU/ALU/_825_ ( .A(\EXU/casez_tmp_0 [7] ), .Z(\EXU/ALU/_164_ ) );
BUF_X1 \EXU/ALU/_826_ ( .A(\EXU/_0029_ ), .Z(\EXU/ALU/_132_ ) );
BUF_X1 \EXU/ALU/_827_ ( .A(\EXU/ALU/_barrelShift_io_out [7] ), .Z(\EXU/ALU/_068_ ) );
BUF_X1 \EXU/ALU/_828_ ( .A(\EXU/ALU/_adder_io_result [7] ), .Z(\EXU/ALU/_031_ ) );
BUF_X1 \EXU/ALU/_829_ ( .A(\EXU/ALU/_100_ ), .Z(\_EXU_io_LSUIn_bits_raddr [7] ) );
BUF_X1 \EXU/ALU/_830_ ( .A(\EXU/casez_tmp_0 [8] ), .Z(\EXU/ALU/_165_ ) );
BUF_X1 \EXU/ALU/_831_ ( .A(\EXU/_0030_ ), .Z(\EXU/ALU/_133_ ) );
BUF_X1 \EXU/ALU/_832_ ( .A(\EXU/ALU/_barrelShift_io_out [8] ), .Z(\EXU/ALU/_069_ ) );
BUF_X1 \EXU/ALU/_833_ ( .A(\EXU/ALU/_adder_io_result [8] ), .Z(\EXU/ALU/_032_ ) );
BUF_X1 \EXU/ALU/_834_ ( .A(\EXU/ALU/_101_ ), .Z(\_EXU_io_LSUIn_bits_raddr [8] ) );
BUF_X1 \EXU/ALU/_835_ ( .A(\EXU/casez_tmp_0 [9] ), .Z(\EXU/ALU/_166_ ) );
BUF_X1 \EXU/ALU/_836_ ( .A(\EXU/_0031_ ), .Z(\EXU/ALU/_134_ ) );
BUF_X1 \EXU/ALU/_837_ ( .A(\EXU/ALU/_barrelShift_io_out [9] ), .Z(\EXU/ALU/_070_ ) );
BUF_X1 \EXU/ALU/_838_ ( .A(\EXU/ALU/_adder_io_result [9] ), .Z(\EXU/ALU/_033_ ) );
BUF_X1 \EXU/ALU/_839_ ( .A(\EXU/ALU/_102_ ), .Z(\_EXU_io_LSUIn_bits_raddr [9] ) );
BUF_X1 \EXU/ALU/_840_ ( .A(\EXU/casez_tmp_0 [10] ), .Z(\EXU/ALU/_136_ ) );
BUF_X1 \EXU/ALU/_841_ ( .A(\EXU/_0001_ ), .Z(\EXU/ALU/_104_ ) );
BUF_X1 \EXU/ALU/_842_ ( .A(\EXU/ALU/_barrelShift_io_out [10] ), .Z(\EXU/ALU/_040_ ) );
BUF_X1 \EXU/ALU/_843_ ( .A(\EXU/ALU/_adder_io_result [10] ), .Z(\EXU/ALU/_003_ ) );
BUF_X1 \EXU/ALU/_844_ ( .A(\EXU/ALU/_072_ ), .Z(\_EXU_io_LSUIn_bits_raddr [10] ) );
BUF_X1 \EXU/ALU/_845_ ( .A(\EXU/casez_tmp_0 [11] ), .Z(\EXU/ALU/_137_ ) );
BUF_X1 \EXU/ALU/_846_ ( .A(\EXU/_0002_ ), .Z(\EXU/ALU/_105_ ) );
BUF_X1 \EXU/ALU/_847_ ( .A(\EXU/ALU/_barrelShift_io_out [11] ), .Z(\EXU/ALU/_041_ ) );
BUF_X1 \EXU/ALU/_848_ ( .A(\EXU/ALU/_adder_io_result [11] ), .Z(\EXU/ALU/_004_ ) );
BUF_X1 \EXU/ALU/_849_ ( .A(\EXU/ALU/_073_ ), .Z(\_EXU_io_LSUIn_bits_raddr [11] ) );
BUF_X1 \EXU/ALU/_850_ ( .A(\EXU/casez_tmp_0 [12] ), .Z(\EXU/ALU/_138_ ) );
BUF_X1 \EXU/ALU/_851_ ( .A(\EXU/_0003_ ), .Z(\EXU/ALU/_106_ ) );
BUF_X1 \EXU/ALU/_852_ ( .A(\EXU/ALU/_barrelShift_io_out [12] ), .Z(\EXU/ALU/_042_ ) );
BUF_X1 \EXU/ALU/_853_ ( .A(\EXU/ALU/_adder_io_result [12] ), .Z(\EXU/ALU/_005_ ) );
BUF_X1 \EXU/ALU/_854_ ( .A(\EXU/ALU/_074_ ), .Z(\_EXU_io_LSUIn_bits_raddr [12] ) );
BUF_X1 \EXU/ALU/_855_ ( .A(\EXU/casez_tmp_0 [13] ), .Z(\EXU/ALU/_139_ ) );
BUF_X1 \EXU/ALU/_856_ ( .A(\EXU/_0004_ ), .Z(\EXU/ALU/_107_ ) );
BUF_X1 \EXU/ALU/_857_ ( .A(\EXU/ALU/_barrelShift_io_out [13] ), .Z(\EXU/ALU/_043_ ) );
BUF_X1 \EXU/ALU/_858_ ( .A(\EXU/ALU/_adder_io_result [13] ), .Z(\EXU/ALU/_006_ ) );
BUF_X1 \EXU/ALU/_859_ ( .A(\EXU/ALU/_075_ ), .Z(\_EXU_io_LSUIn_bits_raddr [13] ) );
BUF_X1 \EXU/ALU/_860_ ( .A(\EXU/casez_tmp_0 [14] ), .Z(\EXU/ALU/_140_ ) );
BUF_X1 \EXU/ALU/_861_ ( .A(\EXU/_0005_ ), .Z(\EXU/ALU/_108_ ) );
BUF_X1 \EXU/ALU/_862_ ( .A(\EXU/ALU/_barrelShift_io_out [14] ), .Z(\EXU/ALU/_044_ ) );
BUF_X1 \EXU/ALU/_863_ ( .A(\EXU/ALU/_adder_io_result [14] ), .Z(\EXU/ALU/_007_ ) );
BUF_X1 \EXU/ALU/_864_ ( .A(\EXU/ALU/_076_ ), .Z(\_EXU_io_LSUIn_bits_raddr [14] ) );
BUF_X1 \EXU/ALU/_865_ ( .A(\EXU/casez_tmp_0 [15] ), .Z(\EXU/ALU/_141_ ) );
BUF_X1 \EXU/ALU/_866_ ( .A(\EXU/_0006_ ), .Z(\EXU/ALU/_109_ ) );
BUF_X1 \EXU/ALU/_867_ ( .A(\EXU/ALU/_barrelShift_io_out [15] ), .Z(\EXU/ALU/_045_ ) );
BUF_X1 \EXU/ALU/_868_ ( .A(\EXU/ALU/_adder_io_result [15] ), .Z(\EXU/ALU/_008_ ) );
BUF_X1 \EXU/ALU/_869_ ( .A(\EXU/ALU/_077_ ), .Z(\_EXU_io_LSUIn_bits_raddr [15] ) );
BUF_X1 \EXU/ALU/_870_ ( .A(\EXU/casez_tmp_0 [16] ), .Z(\EXU/ALU/_142_ ) );
BUF_X1 \EXU/ALU/_871_ ( .A(\EXU/_0007_ ), .Z(\EXU/ALU/_110_ ) );
BUF_X1 \EXU/ALU/_872_ ( .A(\EXU/ALU/_barrelShift_io_out [16] ), .Z(\EXU/ALU/_046_ ) );
BUF_X1 \EXU/ALU/_873_ ( .A(\EXU/ALU/_adder_io_result [16] ), .Z(\EXU/ALU/_009_ ) );
BUF_X1 \EXU/ALU/_874_ ( .A(\EXU/ALU/_078_ ), .Z(\_EXU_io_LSUIn_bits_raddr [16] ) );
BUF_X1 \EXU/ALU/_875_ ( .A(\EXU/casez_tmp_0 [17] ), .Z(\EXU/ALU/_143_ ) );
BUF_X1 \EXU/ALU/_876_ ( .A(\EXU/_0008_ ), .Z(\EXU/ALU/_111_ ) );
BUF_X1 \EXU/ALU/_877_ ( .A(\EXU/ALU/_barrelShift_io_out [17] ), .Z(\EXU/ALU/_047_ ) );
BUF_X1 \EXU/ALU/_878_ ( .A(\EXU/ALU/_adder_io_result [17] ), .Z(\EXU/ALU/_010_ ) );
BUF_X1 \EXU/ALU/_879_ ( .A(\EXU/ALU/_079_ ), .Z(\_EXU_io_LSUIn_bits_raddr [17] ) );
BUF_X1 \EXU/ALU/_880_ ( .A(\EXU/casez_tmp_0 [18] ), .Z(\EXU/ALU/_144_ ) );
BUF_X1 \EXU/ALU/_881_ ( .A(\EXU/_0009_ ), .Z(\EXU/ALU/_112_ ) );
BUF_X1 \EXU/ALU/_882_ ( .A(\EXU/ALU/_barrelShift_io_out [18] ), .Z(\EXU/ALU/_048_ ) );
BUF_X1 \EXU/ALU/_883_ ( .A(\EXU/ALU/_adder_io_result [18] ), .Z(\EXU/ALU/_011_ ) );
BUF_X1 \EXU/ALU/_884_ ( .A(\EXU/ALU/_080_ ), .Z(\_EXU_io_LSUIn_bits_raddr [18] ) );
BUF_X1 \EXU/ALU/_885_ ( .A(\EXU/casez_tmp_0 [19] ), .Z(\EXU/ALU/_145_ ) );
BUF_X1 \EXU/ALU/_886_ ( .A(\EXU/_0010_ ), .Z(\EXU/ALU/_113_ ) );
BUF_X1 \EXU/ALU/_887_ ( .A(\EXU/ALU/_barrelShift_io_out [19] ), .Z(\EXU/ALU/_049_ ) );
BUF_X1 \EXU/ALU/_888_ ( .A(\EXU/ALU/_adder_io_result [19] ), .Z(\EXU/ALU/_012_ ) );
BUF_X1 \EXU/ALU/_889_ ( .A(\EXU/ALU/_081_ ), .Z(\_EXU_io_LSUIn_bits_raddr [19] ) );
BUF_X1 \EXU/ALU/_890_ ( .A(\EXU/casez_tmp_0 [20] ), .Z(\EXU/ALU/_147_ ) );
BUF_X1 \EXU/ALU/_891_ ( .A(\EXU/_0012_ ), .Z(\EXU/ALU/_115_ ) );
BUF_X1 \EXU/ALU/_892_ ( .A(\EXU/ALU/_barrelShift_io_out [20] ), .Z(\EXU/ALU/_051_ ) );
BUF_X1 \EXU/ALU/_893_ ( .A(\EXU/ALU/_adder_io_result [20] ), .Z(\EXU/ALU/_014_ ) );
BUF_X1 \EXU/ALU/_894_ ( .A(\EXU/ALU/_083_ ), .Z(\_EXU_io_LSUIn_bits_raddr [20] ) );
BUF_X1 \EXU/ALU/_895_ ( .A(\EXU/casez_tmp_0 [21] ), .Z(\EXU/ALU/_148_ ) );
BUF_X1 \EXU/ALU/_896_ ( .A(\EXU/_0013_ ), .Z(\EXU/ALU/_116_ ) );
BUF_X1 \EXU/ALU/_897_ ( .A(\EXU/ALU/_barrelShift_io_out [21] ), .Z(\EXU/ALU/_052_ ) );
BUF_X1 \EXU/ALU/_898_ ( .A(\EXU/ALU/_adder_io_result [21] ), .Z(\EXU/ALU/_015_ ) );
BUF_X1 \EXU/ALU/_899_ ( .A(\EXU/ALU/_084_ ), .Z(\_EXU_io_LSUIn_bits_raddr [21] ) );
BUF_X1 \EXU/ALU/_900_ ( .A(\EXU/casez_tmp_0 [22] ), .Z(\EXU/ALU/_149_ ) );
BUF_X1 \EXU/ALU/_901_ ( .A(\EXU/_0014_ ), .Z(\EXU/ALU/_117_ ) );
BUF_X1 \EXU/ALU/_902_ ( .A(\EXU/ALU/_barrelShift_io_out [22] ), .Z(\EXU/ALU/_053_ ) );
BUF_X1 \EXU/ALU/_903_ ( .A(\EXU/ALU/_adder_io_result [22] ), .Z(\EXU/ALU/_016_ ) );
BUF_X1 \EXU/ALU/_904_ ( .A(\EXU/ALU/_085_ ), .Z(\_EXU_io_LSUIn_bits_raddr [22] ) );
BUF_X1 \EXU/ALU/_905_ ( .A(\EXU/casez_tmp_0 [23] ), .Z(\EXU/ALU/_150_ ) );
BUF_X1 \EXU/ALU/_906_ ( .A(\EXU/_0015_ ), .Z(\EXU/ALU/_118_ ) );
BUF_X1 \EXU/ALU/_907_ ( .A(\EXU/ALU/_barrelShift_io_out [23] ), .Z(\EXU/ALU/_054_ ) );
BUF_X1 \EXU/ALU/_908_ ( .A(\EXU/ALU/_adder_io_result [23] ), .Z(\EXU/ALU/_017_ ) );
BUF_X1 \EXU/ALU/_909_ ( .A(\EXU/ALU/_086_ ), .Z(\_EXU_io_LSUIn_bits_raddr [23] ) );
BUF_X1 \EXU/ALU/_910_ ( .A(\EXU/casez_tmp_0 [24] ), .Z(\EXU/ALU/_151_ ) );
BUF_X1 \EXU/ALU/_911_ ( .A(\EXU/_0016_ ), .Z(\EXU/ALU/_119_ ) );
BUF_X1 \EXU/ALU/_912_ ( .A(\EXU/ALU/_barrelShift_io_out [24] ), .Z(\EXU/ALU/_055_ ) );
BUF_X1 \EXU/ALU/_913_ ( .A(\EXU/ALU/_adder_io_result [24] ), .Z(\EXU/ALU/_018_ ) );
BUF_X1 \EXU/ALU/_914_ ( .A(\EXU/ALU/_087_ ), .Z(\_EXU_io_LSUIn_bits_raddr [24] ) );
BUF_X1 \EXU/ALU/_915_ ( .A(\EXU/casez_tmp_0 [25] ), .Z(\EXU/ALU/_152_ ) );
BUF_X1 \EXU/ALU/_916_ ( .A(\EXU/_0017_ ), .Z(\EXU/ALU/_120_ ) );
BUF_X1 \EXU/ALU/_917_ ( .A(\EXU/ALU/_barrelShift_io_out [25] ), .Z(\EXU/ALU/_056_ ) );
BUF_X1 \EXU/ALU/_918_ ( .A(\EXU/ALU/_adder_io_result [25] ), .Z(\EXU/ALU/_019_ ) );
BUF_X1 \EXU/ALU/_919_ ( .A(\EXU/ALU/_088_ ), .Z(\_EXU_io_LSUIn_bits_raddr [25] ) );
BUF_X1 \EXU/ALU/_920_ ( .A(\EXU/casez_tmp_0 [26] ), .Z(\EXU/ALU/_153_ ) );
BUF_X1 \EXU/ALU/_921_ ( .A(\EXU/_0018_ ), .Z(\EXU/ALU/_121_ ) );
BUF_X1 \EXU/ALU/_922_ ( .A(\EXU/ALU/_barrelShift_io_out [26] ), .Z(\EXU/ALU/_057_ ) );
BUF_X1 \EXU/ALU/_923_ ( .A(\EXU/ALU/_adder_io_result [26] ), .Z(\EXU/ALU/_020_ ) );
BUF_X1 \EXU/ALU/_924_ ( .A(\EXU/ALU/_089_ ), .Z(\_EXU_io_LSUIn_bits_raddr [26] ) );
BUF_X1 \EXU/ALU/_925_ ( .A(\EXU/casez_tmp_0 [27] ), .Z(\EXU/ALU/_154_ ) );
BUF_X1 \EXU/ALU/_926_ ( .A(\EXU/_0019_ ), .Z(\EXU/ALU/_122_ ) );
BUF_X1 \EXU/ALU/_927_ ( .A(\EXU/ALU/_barrelShift_io_out [27] ), .Z(\EXU/ALU/_058_ ) );
BUF_X1 \EXU/ALU/_928_ ( .A(\EXU/ALU/_adder_io_result [27] ), .Z(\EXU/ALU/_021_ ) );
BUF_X1 \EXU/ALU/_929_ ( .A(\EXU/ALU/_090_ ), .Z(\_EXU_io_LSUIn_bits_raddr [27] ) );
BUF_X1 \EXU/ALU/_930_ ( .A(\EXU/casez_tmp_0 [28] ), .Z(\EXU/ALU/_155_ ) );
BUF_X1 \EXU/ALU/_931_ ( .A(\EXU/_0020_ ), .Z(\EXU/ALU/_123_ ) );
BUF_X1 \EXU/ALU/_932_ ( .A(\EXU/ALU/_barrelShift_io_out [28] ), .Z(\EXU/ALU/_059_ ) );
BUF_X1 \EXU/ALU/_933_ ( .A(\EXU/ALU/_adder_io_result [28] ), .Z(\EXU/ALU/_022_ ) );
BUF_X1 \EXU/ALU/_934_ ( .A(\EXU/ALU/_091_ ), .Z(\_EXU_io_LSUIn_bits_raddr [28] ) );
BUF_X1 \EXU/ALU/_935_ ( .A(\EXU/casez_tmp_0 [29] ), .Z(\EXU/ALU/_156_ ) );
BUF_X1 \EXU/ALU/_936_ ( .A(\EXU/_0021_ ), .Z(\EXU/ALU/_124_ ) );
BUF_X1 \EXU/ALU/_937_ ( .A(\EXU/ALU/_barrelShift_io_out [29] ), .Z(\EXU/ALU/_060_ ) );
BUF_X1 \EXU/ALU/_938_ ( .A(\EXU/ALU/_adder_io_result [29] ), .Z(\EXU/ALU/_023_ ) );
BUF_X1 \EXU/ALU/_939_ ( .A(\EXU/ALU/_092_ ), .Z(\_EXU_io_LSUIn_bits_raddr [29] ) );
BUF_X1 \EXU/ALU/_940_ ( .A(\EXU/casez_tmp_0 [30] ), .Z(\EXU/ALU/_158_ ) );
BUF_X1 \EXU/ALU/_941_ ( .A(\EXU/_0023_ ), .Z(\EXU/ALU/_126_ ) );
BUF_X1 \EXU/ALU/_942_ ( .A(\EXU/ALU/_barrelShift_io_out [30] ), .Z(\EXU/ALU/_062_ ) );
BUF_X1 \EXU/ALU/_943_ ( .A(\EXU/ALU/_adder_io_result [30] ), .Z(\EXU/ALU/_025_ ) );
BUF_X1 \EXU/ALU/_944_ ( .A(\EXU/ALU/_094_ ), .Z(\_EXU_io_LSUIn_bits_raddr [30] ) );
BUF_X1 \EXU/ALU/_945_ ( .A(\EXU/casez_tmp_0 [31] ), .Z(\EXU/ALU/_159_ ) );
BUF_X1 \EXU/ALU/_946_ ( .A(\EXU/_0024_ ), .Z(\EXU/ALU/_127_ ) );
BUF_X1 \EXU/ALU/_947_ ( .A(\EXU/ALU/_barrelShift_io_out [31] ), .Z(\EXU/ALU/_063_ ) );
BUF_X1 \EXU/ALU/_948_ ( .A(\EXU/ALU/_095_ ), .Z(\_EXU_io_LSUIn_bits_raddr [31] ) );
XOR2_X1 \EXU/ALU/adder/_371_ ( .A(\EXU/ALU/adder/_034_ ), .B(\EXU/ALU/adder/_002_ ), .Z(\EXU/ALU/adder/_067_ ) );
XNOR2_X2 \EXU/ALU/adder/_372_ ( .A(fanout_net_16 ), .B(\EXU/ALU/adder/_045_ ), .ZN(\EXU/ALU/adder/_100_ ) );
XNOR2_X1 \EXU/ALU/adder/_373_ ( .A(\EXU/ALU/adder/_100_ ), .B(\EXU/ALU/adder/_013_ ), .ZN(\EXU/ALU/adder/_101_ ) );
INV_X1 \EXU/ALU/adder/_374_ ( .A(\EXU/ALU/adder/_034_ ), .ZN(\EXU/ALU/adder/_102_ ) );
NOR2_X1 \EXU/ALU/adder/_375_ ( .A1(\EXU/ALU/adder/_102_ ), .A2(\EXU/ALU/adder/_002_ ), .ZN(\EXU/ALU/adder/_103_ ) );
NOR2_X1 \EXU/ALU/adder/_376_ ( .A1(\EXU/ALU/adder/_034_ ), .A2(fanout_net_16 ), .ZN(\EXU/ALU/adder/_104_ ) );
NOR2_X1 \EXU/ALU/adder/_377_ ( .A1(\EXU/ALU/adder/_103_ ), .A2(\EXU/ALU/adder/_104_ ), .ZN(\EXU/ALU/adder/_105_ ) );
XOR2_X1 \EXU/ALU/adder/_378_ ( .A(\EXU/ALU/adder/_101_ ), .B(\EXU/ALU/adder/_105_ ), .Z(\EXU/ALU/adder/_078_ ) );
NAND2_X1 \EXU/ALU/adder/_379_ ( .A1(\EXU/ALU/adder/_101_ ), .A2(\EXU/ALU/adder/_105_ ), .ZN(\EXU/ALU/adder/_106_ ) );
INV_X1 \EXU/ALU/adder/_380_ ( .A(\EXU/ALU/adder/_013_ ), .ZN(\EXU/ALU/adder/_107_ ) );
OR2_X1 \EXU/ALU/adder/_381_ ( .A1(\EXU/ALU/adder/_100_ ), .A2(\EXU/ALU/adder/_107_ ), .ZN(\EXU/ALU/adder/_108_ ) );
XNOR2_X2 \EXU/ALU/adder/_382_ ( .A(fanout_net_16 ), .B(\EXU/ALU/adder/_056_ ), .ZN(\EXU/ALU/adder/_109_ ) );
INV_X1 \EXU/ALU/adder/_383_ ( .A(\EXU/ALU/adder/_024_ ), .ZN(\EXU/ALU/adder/_110_ ) );
XNOR2_X1 \EXU/ALU/adder/_384_ ( .A(\EXU/ALU/adder/_109_ ), .B(\EXU/ALU/adder/_110_ ), .ZN(\EXU/ALU/adder/_111_ ) );
AND3_X1 \EXU/ALU/adder/_385_ ( .A1(\EXU/ALU/adder/_106_ ), .A2(\EXU/ALU/adder/_108_ ), .A3(\EXU/ALU/adder/_111_ ), .ZN(\EXU/ALU/adder/_112_ ) );
AOI21_X2 \EXU/ALU/adder/_386_ ( .A(\EXU/ALU/adder/_111_ ), .B1(\EXU/ALU/adder/_106_ ), .B2(\EXU/ALU/adder/_108_ ), .ZN(\EXU/ALU/adder/_113_ ) );
NOR2_X1 \EXU/ALU/adder/_387_ ( .A1(\EXU/ALU/adder/_112_ ), .A2(\EXU/ALU/adder/_113_ ), .ZN(\EXU/ALU/adder/_089_ ) );
NOR2_X1 \EXU/ALU/adder/_388_ ( .A1(\EXU/ALU/adder/_109_ ), .A2(\EXU/ALU/adder/_110_ ), .ZN(\EXU/ALU/adder/_114_ ) );
NOR2_X1 \EXU/ALU/adder/_389_ ( .A1(\EXU/ALU/adder/_113_ ), .A2(\EXU/ALU/adder/_114_ ), .ZN(\EXU/ALU/adder/_115_ ) );
XNOR2_X2 \EXU/ALU/adder/_390_ ( .A(fanout_net_16 ), .B(\EXU/ALU/adder/_059_ ), .ZN(\EXU/ALU/adder/_116_ ) );
INV_X1 \EXU/ALU/adder/_391_ ( .A(\EXU/ALU/adder/_027_ ), .ZN(\EXU/ALU/adder/_117_ ) );
XNOR2_X2 \EXU/ALU/adder/_392_ ( .A(\EXU/ALU/adder/_116_ ), .B(\EXU/ALU/adder/_117_ ), .ZN(\EXU/ALU/adder/_118_ ) );
XNOR2_X1 \EXU/ALU/adder/_393_ ( .A(\EXU/ALU/adder/_115_ ), .B(\EXU/ALU/adder/_118_ ), .ZN(\EXU/ALU/adder/_119_ ) );
INV_X1 \EXU/ALU/adder/_394_ ( .A(\EXU/ALU/adder/_119_ ), .ZN(\EXU/ALU/adder/_092_ ) );
AOI211_X2 \EXU/ALU/adder/_395_ ( .A(\EXU/ALU/adder/_111_ ), .B(\EXU/ALU/adder/_118_ ), .C1(\EXU/ALU/adder/_106_ ), .C2(\EXU/ALU/adder/_108_ ), .ZN(\EXU/ALU/adder/_120_ ) );
OR3_X4 \EXU/ALU/adder/_396_ ( .A1(\EXU/ALU/adder/_118_ ), .A2(\EXU/ALU/adder/_110_ ), .A3(\EXU/ALU/adder/_109_ ), .ZN(\EXU/ALU/adder/_121_ ) );
OAI21_X1 \EXU/ALU/adder/_397_ ( .A(\EXU/ALU/adder/_121_ ), .B1(\EXU/ALU/adder/_117_ ), .B2(\EXU/ALU/adder/_116_ ), .ZN(\EXU/ALU/adder/_122_ ) );
NOR2_X2 \EXU/ALU/adder/_398_ ( .A1(\EXU/ALU/adder/_120_ ), .A2(\EXU/ALU/adder/_122_ ), .ZN(\EXU/ALU/adder/_123_ ) );
XNOR2_X2 \EXU/ALU/adder/_399_ ( .A(fanout_net_16 ), .B(\EXU/ALU/adder/_060_ ), .ZN(\EXU/ALU/adder/_124_ ) );
XNOR2_X1 \EXU/ALU/adder/_400_ ( .A(\EXU/ALU/adder/_124_ ), .B(\EXU/ALU/adder/_028_ ), .ZN(\EXU/ALU/adder/_125_ ) );
XNOR2_X1 \EXU/ALU/adder/_401_ ( .A(\EXU/ALU/adder/_123_ ), .B(\EXU/ALU/adder/_125_ ), .ZN(\EXU/ALU/adder/_093_ ) );
INV_X1 \EXU/ALU/adder/_402_ ( .A(\EXU/ALU/adder/_028_ ), .ZN(\EXU/ALU/adder/_126_ ) );
NOR2_X2 \EXU/ALU/adder/_403_ ( .A1(\EXU/ALU/adder/_124_ ), .A2(\EXU/ALU/adder/_126_ ), .ZN(\EXU/ALU/adder/_127_ ) );
AND2_X1 \EXU/ALU/adder/_404_ ( .A1(\EXU/ALU/adder/_124_ ), .A2(\EXU/ALU/adder/_126_ ), .ZN(\EXU/ALU/adder/_128_ ) );
NOR3_X1 \EXU/ALU/adder/_405_ ( .A1(\EXU/ALU/adder/_123_ ), .A2(\EXU/ALU/adder/_127_ ), .A3(\EXU/ALU/adder/_128_ ), .ZN(\EXU/ALU/adder/_129_ ) );
NOR2_X1 \EXU/ALU/adder/_406_ ( .A1(\EXU/ALU/adder/_129_ ), .A2(\EXU/ALU/adder/_127_ ), .ZN(\EXU/ALU/adder/_130_ ) );
XNOR2_X2 \EXU/ALU/adder/_407_ ( .A(fanout_net_16 ), .B(\EXU/ALU/adder/_061_ ), .ZN(\EXU/ALU/adder/_131_ ) );
XNOR2_X2 \EXU/ALU/adder/_408_ ( .A(\EXU/ALU/adder/_131_ ), .B(\EXU/ALU/adder/_029_ ), .ZN(\EXU/ALU/adder/_132_ ) );
INV_X1 \EXU/ALU/adder/_409_ ( .A(\EXU/ALU/adder/_132_ ), .ZN(\EXU/ALU/adder/_133_ ) );
XNOR2_X1 \EXU/ALU/adder/_410_ ( .A(\EXU/ALU/adder/_130_ ), .B(\EXU/ALU/adder/_133_ ), .ZN(\EXU/ALU/adder/_134_ ) );
INV_X1 \EXU/ALU/adder/_411_ ( .A(\EXU/ALU/adder/_134_ ), .ZN(\EXU/ALU/adder/_094_ ) );
NOR4_X1 \EXU/ALU/adder/_412_ ( .A1(\EXU/ALU/adder/_123_ ), .A2(\EXU/ALU/adder/_127_ ), .A3(\EXU/ALU/adder/_128_ ), .A4(\EXU/ALU/adder/_133_ ), .ZN(\EXU/ALU/adder/_135_ ) );
NAND2_X2 \EXU/ALU/adder/_413_ ( .A1(\EXU/ALU/adder/_132_ ), .A2(\EXU/ALU/adder/_127_ ), .ZN(\EXU/ALU/adder/_136_ ) );
INV_X1 \EXU/ALU/adder/_414_ ( .A(\EXU/ALU/adder/_029_ ), .ZN(\EXU/ALU/adder/_137_ ) );
OAI21_X1 \EXU/ALU/adder/_415_ ( .A(\EXU/ALU/adder/_136_ ), .B1(\EXU/ALU/adder/_137_ ), .B2(\EXU/ALU/adder/_131_ ), .ZN(\EXU/ALU/adder/_138_ ) );
OR2_X1 \EXU/ALU/adder/_416_ ( .A1(\EXU/ALU/adder/_135_ ), .A2(\EXU/ALU/adder/_138_ ), .ZN(\EXU/ALU/adder/_139_ ) );
XNOR2_X1 \EXU/ALU/adder/_417_ ( .A(fanout_net_16 ), .B(\EXU/ALU/adder/_062_ ), .ZN(\EXU/ALU/adder/_140_ ) );
XNOR2_X1 \EXU/ALU/adder/_418_ ( .A(\EXU/ALU/adder/_140_ ), .B(\EXU/ALU/adder/_030_ ), .ZN(\EXU/ALU/adder/_141_ ) );
XOR2_X1 \EXU/ALU/adder/_419_ ( .A(\EXU/ALU/adder/_139_ ), .B(\EXU/ALU/adder/_141_ ), .Z(\EXU/ALU/adder/_095_ ) );
AND2_X1 \EXU/ALU/adder/_420_ ( .A1(\EXU/ALU/adder/_139_ ), .A2(\EXU/ALU/adder/_141_ ), .ZN(\EXU/ALU/adder/_142_ ) );
INV_X1 \EXU/ALU/adder/_421_ ( .A(\EXU/ALU/adder/_030_ ), .ZN(\EXU/ALU/adder/_143_ ) );
NOR2_X1 \EXU/ALU/adder/_422_ ( .A1(\EXU/ALU/adder/_140_ ), .A2(\EXU/ALU/adder/_143_ ), .ZN(\EXU/ALU/adder/_144_ ) );
NOR2_X1 \EXU/ALU/adder/_423_ ( .A1(\EXU/ALU/adder/_142_ ), .A2(\EXU/ALU/adder/_144_ ), .ZN(\EXU/ALU/adder/_145_ ) );
XNOR2_X2 \EXU/ALU/adder/_424_ ( .A(fanout_net_16 ), .B(\EXU/ALU/adder/_063_ ), .ZN(\EXU/ALU/adder/_146_ ) );
XNOR2_X2 \EXU/ALU/adder/_425_ ( .A(\EXU/ALU/adder/_146_ ), .B(\EXU/ALU/adder/_031_ ), .ZN(\EXU/ALU/adder/_147_ ) );
XNOR2_X1 \EXU/ALU/adder/_426_ ( .A(\EXU/ALU/adder/_145_ ), .B(\EXU/ALU/adder/_147_ ), .ZN(\EXU/ALU/adder/_096_ ) );
XNOR2_X1 \EXU/ALU/adder/_427_ ( .A(fanout_net_16 ), .B(\EXU/ALU/adder/_064_ ), .ZN(\EXU/ALU/adder/_148_ ) );
XNOR2_X1 \EXU/ALU/adder/_428_ ( .A(\EXU/ALU/adder/_148_ ), .B(\EXU/ALU/adder/_032_ ), .ZN(\EXU/ALU/adder/_149_ ) );
INV_X1 \EXU/ALU/adder/_429_ ( .A(\EXU/ALU/adder/_031_ ), .ZN(\EXU/ALU/adder/_150_ ) );
NOR2_X1 \EXU/ALU/adder/_430_ ( .A1(\EXU/ALU/adder/_146_ ), .A2(\EXU/ALU/adder/_150_ ), .ZN(\EXU/ALU/adder/_151_ ) );
AND3_X2 \EXU/ALU/adder/_431_ ( .A1(\EXU/ALU/adder/_138_ ), .A2(\EXU/ALU/adder/_141_ ), .A3(\EXU/ALU/adder/_147_ ), .ZN(\EXU/ALU/adder/_152_ ) );
AOI211_X2 \EXU/ALU/adder/_432_ ( .A(\EXU/ALU/adder/_151_ ), .B(\EXU/ALU/adder/_152_ ), .C1(\EXU/ALU/adder/_144_ ), .C2(\EXU/ALU/adder/_147_ ), .ZN(\EXU/ALU/adder/_153_ ) );
INV_X2 \EXU/ALU/adder/_433_ ( .A(\EXU/ALU/adder/_153_ ), .ZN(\EXU/ALU/adder/_154_ ) );
NAND4_X1 \EXU/ALU/adder/_434_ ( .A1(\EXU/ALU/adder/_125_ ), .A2(\EXU/ALU/adder/_132_ ), .A3(\EXU/ALU/adder/_141_ ), .A4(\EXU/ALU/adder/_147_ ), .ZN(\EXU/ALU/adder/_155_ ) );
NOR2_X4 \EXU/ALU/adder/_435_ ( .A1(\EXU/ALU/adder/_123_ ), .A2(\EXU/ALU/adder/_155_ ), .ZN(\EXU/ALU/adder/_156_ ) );
OAI21_X1 \EXU/ALU/adder/_436_ ( .A(\EXU/ALU/adder/_149_ ), .B1(\EXU/ALU/adder/_154_ ), .B2(\EXU/ALU/adder/_156_ ), .ZN(\EXU/ALU/adder/_157_ ) );
OR3_X2 \EXU/ALU/adder/_437_ ( .A1(\EXU/ALU/adder/_154_ ), .A2(\EXU/ALU/adder/_156_ ), .A3(\EXU/ALU/adder/_149_ ), .ZN(\EXU/ALU/adder/_158_ ) );
AND2_X2 \EXU/ALU/adder/_438_ ( .A1(\EXU/ALU/adder/_157_ ), .A2(\EXU/ALU/adder/_158_ ), .ZN(\EXU/ALU/adder/_097_ ) );
INV_X1 \EXU/ALU/adder/_439_ ( .A(\EXU/ALU/adder/_032_ ), .ZN(\EXU/ALU/adder/_159_ ) );
NOR2_X1 \EXU/ALU/adder/_440_ ( .A1(\EXU/ALU/adder/_148_ ), .A2(\EXU/ALU/adder/_159_ ), .ZN(\EXU/ALU/adder/_160_ ) );
INV_X1 \EXU/ALU/adder/_441_ ( .A(\EXU/ALU/adder/_160_ ), .ZN(\EXU/ALU/adder/_161_ ) );
AND2_X1 \EXU/ALU/adder/_442_ ( .A1(\EXU/ALU/adder/_157_ ), .A2(\EXU/ALU/adder/_161_ ), .ZN(\EXU/ALU/adder/_162_ ) );
XNOR2_X2 \EXU/ALU/adder/_443_ ( .A(fanout_net_16 ), .B(\EXU/ALU/adder/_065_ ), .ZN(\EXU/ALU/adder/_163_ ) );
XNOR2_X2 \EXU/ALU/adder/_444_ ( .A(\EXU/ALU/adder/_163_ ), .B(\EXU/ALU/adder/_033_ ), .ZN(\EXU/ALU/adder/_164_ ) );
XNOR2_X1 \EXU/ALU/adder/_445_ ( .A(\EXU/ALU/adder/_162_ ), .B(\EXU/ALU/adder/_164_ ), .ZN(\EXU/ALU/adder/_098_ ) );
XNOR2_X1 \EXU/ALU/adder/_446_ ( .A(fanout_net_16 ), .B(\EXU/ALU/adder/_035_ ), .ZN(\EXU/ALU/adder/_165_ ) );
XNOR2_X1 \EXU/ALU/adder/_447_ ( .A(\EXU/ALU/adder/_165_ ), .B(\EXU/ALU/adder/_003_ ), .ZN(\EXU/ALU/adder/_166_ ) );
NAND2_X1 \EXU/ALU/adder/_448_ ( .A1(\EXU/ALU/adder/_164_ ), .A2(\EXU/ALU/adder/_149_ ), .ZN(\EXU/ALU/adder/_167_ ) );
INV_X1 \EXU/ALU/adder/_449_ ( .A(\EXU/ALU/adder/_156_ ), .ZN(\EXU/ALU/adder/_168_ ) );
AOI21_X1 \EXU/ALU/adder/_450_ ( .A(\EXU/ALU/adder/_167_ ), .B1(\EXU/ALU/adder/_168_ ), .B2(\EXU/ALU/adder/_153_ ), .ZN(\EXU/ALU/adder/_169_ ) );
NAND2_X1 \EXU/ALU/adder/_451_ ( .A1(\EXU/ALU/adder/_164_ ), .A2(\EXU/ALU/adder/_160_ ), .ZN(\EXU/ALU/adder/_170_ ) );
INV_X1 \EXU/ALU/adder/_452_ ( .A(\EXU/ALU/adder/_033_ ), .ZN(\EXU/ALU/adder/_171_ ) );
OAI21_X1 \EXU/ALU/adder/_453_ ( .A(\EXU/ALU/adder/_170_ ), .B1(\EXU/ALU/adder/_171_ ), .B2(\EXU/ALU/adder/_163_ ), .ZN(\EXU/ALU/adder/_172_ ) );
OAI21_X1 \EXU/ALU/adder/_454_ ( .A(\EXU/ALU/adder/_166_ ), .B1(\EXU/ALU/adder/_169_ ), .B2(\EXU/ALU/adder/_172_ ), .ZN(\EXU/ALU/adder/_173_ ) );
OR3_X2 \EXU/ALU/adder/_455_ ( .A1(\EXU/ALU/adder/_169_ ), .A2(\EXU/ALU/adder/_172_ ), .A3(\EXU/ALU/adder/_166_ ), .ZN(\EXU/ALU/adder/_174_ ) );
AND2_X1 \EXU/ALU/adder/_456_ ( .A1(\EXU/ALU/adder/_173_ ), .A2(\EXU/ALU/adder/_174_ ), .ZN(\EXU/ALU/adder/_068_ ) );
INV_X1 \EXU/ALU/adder/_457_ ( .A(\EXU/ALU/adder/_003_ ), .ZN(\EXU/ALU/adder/_175_ ) );
NOR2_X1 \EXU/ALU/adder/_458_ ( .A1(\EXU/ALU/adder/_165_ ), .A2(\EXU/ALU/adder/_175_ ), .ZN(\EXU/ALU/adder/_176_ ) );
INV_X1 \EXU/ALU/adder/_459_ ( .A(\EXU/ALU/adder/_176_ ), .ZN(\EXU/ALU/adder/_177_ ) );
NAND2_X1 \EXU/ALU/adder/_460_ ( .A1(\EXU/ALU/adder/_173_ ), .A2(\EXU/ALU/adder/_177_ ), .ZN(\EXU/ALU/adder/_178_ ) );
XNOR2_X2 \EXU/ALU/adder/_461_ ( .A(fanout_net_16 ), .B(\EXU/ALU/adder/_036_ ), .ZN(\EXU/ALU/adder/_179_ ) );
XNOR2_X2 \EXU/ALU/adder/_462_ ( .A(\EXU/ALU/adder/_179_ ), .B(\EXU/ALU/adder/_004_ ), .ZN(\EXU/ALU/adder/_180_ ) );
XNOR2_X1 \EXU/ALU/adder/_463_ ( .A(\EXU/ALU/adder/_178_ ), .B(\EXU/ALU/adder/_180_ ), .ZN(\EXU/ALU/adder/_181_ ) );
INV_X1 \EXU/ALU/adder/_464_ ( .A(\EXU/ALU/adder/_181_ ), .ZN(\EXU/ALU/adder/_069_ ) );
AND2_X1 \EXU/ALU/adder/_465_ ( .A1(\EXU/ALU/adder/_166_ ), .A2(\EXU/ALU/adder/_180_ ), .ZN(\EXU/ALU/adder/_182_ ) );
AND3_X1 \EXU/ALU/adder/_466_ ( .A1(\EXU/ALU/adder/_182_ ), .A2(\EXU/ALU/adder/_149_ ), .A3(\EXU/ALU/adder/_164_ ), .ZN(\EXU/ALU/adder/_183_ ) );
OAI21_X2 \EXU/ALU/adder/_467_ ( .A(\EXU/ALU/adder/_183_ ), .B1(\EXU/ALU/adder/_154_ ), .B2(\EXU/ALU/adder/_156_ ), .ZN(\EXU/ALU/adder/_184_ ) );
NAND2_X1 \EXU/ALU/adder/_468_ ( .A1(\EXU/ALU/adder/_180_ ), .A2(\EXU/ALU/adder/_176_ ), .ZN(\EXU/ALU/adder/_185_ ) );
INV_X1 \EXU/ALU/adder/_469_ ( .A(\EXU/ALU/adder/_004_ ), .ZN(\EXU/ALU/adder/_186_ ) );
OAI21_X1 \EXU/ALU/adder/_470_ ( .A(\EXU/ALU/adder/_185_ ), .B1(\EXU/ALU/adder/_186_ ), .B2(\EXU/ALU/adder/_179_ ), .ZN(\EXU/ALU/adder/_187_ ) );
AOI21_X2 \EXU/ALU/adder/_471_ ( .A(\EXU/ALU/adder/_187_ ), .B1(\EXU/ALU/adder/_172_ ), .B2(\EXU/ALU/adder/_182_ ), .ZN(\EXU/ALU/adder/_188_ ) );
AND2_X2 \EXU/ALU/adder/_472_ ( .A1(\EXU/ALU/adder/_184_ ), .A2(\EXU/ALU/adder/_188_ ), .ZN(\EXU/ALU/adder/_189_ ) );
XNOR2_X1 \EXU/ALU/adder/_473_ ( .A(fanout_net_16 ), .B(\EXU/ALU/adder/_037_ ), .ZN(\EXU/ALU/adder/_190_ ) );
XNOR2_X1 \EXU/ALU/adder/_474_ ( .A(\EXU/ALU/adder/_190_ ), .B(\EXU/ALU/adder/_005_ ), .ZN(\EXU/ALU/adder/_191_ ) );
XNOR2_X1 \EXU/ALU/adder/_475_ ( .A(\EXU/ALU/adder/_189_ ), .B(\EXU/ALU/adder/_191_ ), .ZN(\EXU/ALU/adder/_070_ ) );
INV_X1 \EXU/ALU/adder/_476_ ( .A(\EXU/ALU/adder/_191_ ), .ZN(\EXU/ALU/adder/_192_ ) );
OR2_X1 \EXU/ALU/adder/_477_ ( .A1(\EXU/ALU/adder/_189_ ), .A2(\EXU/ALU/adder/_192_ ), .ZN(\EXU/ALU/adder/_193_ ) );
INV_X1 \EXU/ALU/adder/_478_ ( .A(\EXU/ALU/adder/_005_ ), .ZN(\EXU/ALU/adder/_194_ ) );
OR2_X1 \EXU/ALU/adder/_479_ ( .A1(\EXU/ALU/adder/_190_ ), .A2(\EXU/ALU/adder/_194_ ), .ZN(\EXU/ALU/adder/_195_ ) );
NAND2_X1 \EXU/ALU/adder/_480_ ( .A1(\EXU/ALU/adder/_193_ ), .A2(\EXU/ALU/adder/_195_ ), .ZN(\EXU/ALU/adder/_196_ ) );
XNOR2_X1 \EXU/ALU/adder/_481_ ( .A(fanout_net_16 ), .B(\EXU/ALU/adder/_038_ ), .ZN(\EXU/ALU/adder/_197_ ) );
XNOR2_X1 \EXU/ALU/adder/_482_ ( .A(\EXU/ALU/adder/_197_ ), .B(\EXU/ALU/adder/_006_ ), .ZN(\EXU/ALU/adder/_198_ ) );
XNOR2_X1 \EXU/ALU/adder/_483_ ( .A(\EXU/ALU/adder/_196_ ), .B(\EXU/ALU/adder/_198_ ), .ZN(\EXU/ALU/adder/_199_ ) );
INV_X1 \EXU/ALU/adder/_484_ ( .A(\EXU/ALU/adder/_199_ ), .ZN(\EXU/ALU/adder/_071_ ) );
INV_X1 \EXU/ALU/adder/_485_ ( .A(\EXU/ALU/adder/_198_ ), .ZN(\EXU/ALU/adder/_200_ ) );
AOI211_X4 \EXU/ALU/adder/_486_ ( .A(\EXU/ALU/adder/_192_ ), .B(\EXU/ALU/adder/_200_ ), .C1(\EXU/ALU/adder/_184_ ), .C2(\EXU/ALU/adder/_188_ ), .ZN(\EXU/ALU/adder/_201_ ) );
OR2_X1 \EXU/ALU/adder/_487_ ( .A1(\EXU/ALU/adder/_200_ ), .A2(\EXU/ALU/adder/_195_ ), .ZN(\EXU/ALU/adder/_202_ ) );
INV_X1 \EXU/ALU/adder/_488_ ( .A(\EXU/ALU/adder/_006_ ), .ZN(\EXU/ALU/adder/_203_ ) );
OAI21_X1 \EXU/ALU/adder/_489_ ( .A(\EXU/ALU/adder/_202_ ), .B1(\EXU/ALU/adder/_203_ ), .B2(\EXU/ALU/adder/_197_ ), .ZN(\EXU/ALU/adder/_204_ ) );
NOR2_X1 \EXU/ALU/adder/_490_ ( .A1(\EXU/ALU/adder/_201_ ), .A2(\EXU/ALU/adder/_204_ ), .ZN(\EXU/ALU/adder/_205_ ) );
XNOR2_X1 \EXU/ALU/adder/_491_ ( .A(fanout_net_16 ), .B(\EXU/ALU/adder/_039_ ), .ZN(\EXU/ALU/adder/_206_ ) );
XNOR2_X1 \EXU/ALU/adder/_492_ ( .A(\EXU/ALU/adder/_206_ ), .B(\EXU/ALU/adder/_007_ ), .ZN(\EXU/ALU/adder/_207_ ) );
XNOR2_X1 \EXU/ALU/adder/_493_ ( .A(\EXU/ALU/adder/_205_ ), .B(\EXU/ALU/adder/_207_ ), .ZN(\EXU/ALU/adder/_072_ ) );
INV_X1 \EXU/ALU/adder/_494_ ( .A(\EXU/ALU/adder/_007_ ), .ZN(\EXU/ALU/adder/_208_ ) );
NOR2_X1 \EXU/ALU/adder/_495_ ( .A1(\EXU/ALU/adder/_206_ ), .A2(\EXU/ALU/adder/_208_ ), .ZN(\EXU/ALU/adder/_209_ ) );
AND2_X1 \EXU/ALU/adder/_496_ ( .A1(\EXU/ALU/adder/_206_ ), .A2(\EXU/ALU/adder/_208_ ), .ZN(\EXU/ALU/adder/_210_ ) );
NOR3_X1 \EXU/ALU/adder/_497_ ( .A1(\EXU/ALU/adder/_205_ ), .A2(\EXU/ALU/adder/_209_ ), .A3(\EXU/ALU/adder/_210_ ), .ZN(\EXU/ALU/adder/_211_ ) );
NOR2_X1 \EXU/ALU/adder/_498_ ( .A1(\EXU/ALU/adder/_211_ ), .A2(\EXU/ALU/adder/_209_ ), .ZN(\EXU/ALU/adder/_212_ ) );
XNOR2_X2 \EXU/ALU/adder/_499_ ( .A(fanout_net_16 ), .B(\EXU/ALU/adder/_040_ ), .ZN(\EXU/ALU/adder/_213_ ) );
XNOR2_X1 \EXU/ALU/adder/_500_ ( .A(\EXU/ALU/adder/_213_ ), .B(\EXU/ALU/adder/_008_ ), .ZN(\EXU/ALU/adder/_214_ ) );
XNOR2_X1 \EXU/ALU/adder/_501_ ( .A(\EXU/ALU/adder/_212_ ), .B(\EXU/ALU/adder/_214_ ), .ZN(\EXU/ALU/adder/_073_ ) );
AND2_X2 \EXU/ALU/adder/_502_ ( .A1(\EXU/ALU/adder/_207_ ), .A2(\EXU/ALU/adder/_214_ ), .ZN(\EXU/ALU/adder/_215_ ) );
AND3_X2 \EXU/ALU/adder/_503_ ( .A1(\EXU/ALU/adder/_215_ ), .A2(\EXU/ALU/adder/_191_ ), .A3(\EXU/ALU/adder/_198_ ), .ZN(\EXU/ALU/adder/_216_ ) );
OAI211_X2 \EXU/ALU/adder/_504_ ( .A(\EXU/ALU/adder/_183_ ), .B(\EXU/ALU/adder/_216_ ), .C1(\EXU/ALU/adder/_154_ ), .C2(\EXU/ALU/adder/_156_ ), .ZN(\EXU/ALU/adder/_217_ ) );
NAND2_X1 \EXU/ALU/adder/_505_ ( .A1(\EXU/ALU/adder/_214_ ), .A2(\EXU/ALU/adder/_209_ ), .ZN(\EXU/ALU/adder/_218_ ) );
INV_X1 \EXU/ALU/adder/_506_ ( .A(\EXU/ALU/adder/_008_ ), .ZN(\EXU/ALU/adder/_219_ ) );
OAI21_X1 \EXU/ALU/adder/_507_ ( .A(\EXU/ALU/adder/_218_ ), .B1(\EXU/ALU/adder/_219_ ), .B2(\EXU/ALU/adder/_213_ ), .ZN(\EXU/ALU/adder/_220_ ) );
INV_X1 \EXU/ALU/adder/_508_ ( .A(\EXU/ALU/adder/_216_ ), .ZN(\EXU/ALU/adder/_221_ ) );
NOR2_X1 \EXU/ALU/adder/_509_ ( .A1(\EXU/ALU/adder/_221_ ), .A2(\EXU/ALU/adder/_188_ ), .ZN(\EXU/ALU/adder/_222_ ) );
AOI211_X2 \EXU/ALU/adder/_510_ ( .A(\EXU/ALU/adder/_220_ ), .B(\EXU/ALU/adder/_222_ ), .C1(\EXU/ALU/adder/_204_ ), .C2(\EXU/ALU/adder/_215_ ), .ZN(\EXU/ALU/adder/_223_ ) );
AND2_X2 \EXU/ALU/adder/_511_ ( .A1(\EXU/ALU/adder/_217_ ), .A2(\EXU/ALU/adder/_223_ ), .ZN(\EXU/ALU/adder/_224_ ) );
XNOR2_X1 \EXU/ALU/adder/_512_ ( .A(fanout_net_16 ), .B(\EXU/ALU/adder/_041_ ), .ZN(\EXU/ALU/adder/_225_ ) );
XNOR2_X1 \EXU/ALU/adder/_513_ ( .A(\EXU/ALU/adder/_225_ ), .B(\EXU/ALU/adder/_009_ ), .ZN(\EXU/ALU/adder/_226_ ) );
XNOR2_X1 \EXU/ALU/adder/_514_ ( .A(\EXU/ALU/adder/_224_ ), .B(\EXU/ALU/adder/_226_ ), .ZN(\EXU/ALU/adder/_074_ ) );
INV_X1 \EXU/ALU/adder/_515_ ( .A(\EXU/ALU/adder/_009_ ), .ZN(\EXU/ALU/adder/_227_ ) );
NOR2_X1 \EXU/ALU/adder/_516_ ( .A1(\EXU/ALU/adder/_225_ ), .A2(\EXU/ALU/adder/_227_ ), .ZN(\EXU/ALU/adder/_228_ ) );
AND2_X1 \EXU/ALU/adder/_517_ ( .A1(\EXU/ALU/adder/_225_ ), .A2(\EXU/ALU/adder/_227_ ), .ZN(\EXU/ALU/adder/_229_ ) );
NOR3_X1 \EXU/ALU/adder/_518_ ( .A1(\EXU/ALU/adder/_224_ ), .A2(\EXU/ALU/adder/_228_ ), .A3(\EXU/ALU/adder/_229_ ), .ZN(\EXU/ALU/adder/_230_ ) );
NOR2_X1 \EXU/ALU/adder/_519_ ( .A1(\EXU/ALU/adder/_230_ ), .A2(\EXU/ALU/adder/_228_ ), .ZN(\EXU/ALU/adder/_231_ ) );
XNOR2_X1 \EXU/ALU/adder/_520_ ( .A(fanout_net_16 ), .B(\EXU/ALU/adder/_042_ ), .ZN(\EXU/ALU/adder/_232_ ) );
XNOR2_X1 \EXU/ALU/adder/_521_ ( .A(\EXU/ALU/adder/_232_ ), .B(\EXU/ALU/adder/_010_ ), .ZN(\EXU/ALU/adder/_233_ ) );
XNOR2_X1 \EXU/ALU/adder/_522_ ( .A(\EXU/ALU/adder/_231_ ), .B(\EXU/ALU/adder/_233_ ), .ZN(\EXU/ALU/adder/_075_ ) );
AND2_X1 \EXU/ALU/adder/_523_ ( .A1(\EXU/ALU/adder/_226_ ), .A2(\EXU/ALU/adder/_233_ ), .ZN(\EXU/ALU/adder/_234_ ) );
INV_X1 \EXU/ALU/adder/_524_ ( .A(\EXU/ALU/adder/_234_ ), .ZN(\EXU/ALU/adder/_235_ ) );
AOI21_X1 \EXU/ALU/adder/_525_ ( .A(\EXU/ALU/adder/_235_ ), .B1(\EXU/ALU/adder/_217_ ), .B2(\EXU/ALU/adder/_223_ ), .ZN(\EXU/ALU/adder/_236_ ) );
NAND2_X1 \EXU/ALU/adder/_526_ ( .A1(\EXU/ALU/adder/_233_ ), .A2(\EXU/ALU/adder/_228_ ), .ZN(\EXU/ALU/adder/_237_ ) );
INV_X1 \EXU/ALU/adder/_527_ ( .A(\EXU/ALU/adder/_010_ ), .ZN(\EXU/ALU/adder/_238_ ) );
OAI21_X1 \EXU/ALU/adder/_528_ ( .A(\EXU/ALU/adder/_237_ ), .B1(\EXU/ALU/adder/_238_ ), .B2(\EXU/ALU/adder/_232_ ), .ZN(\EXU/ALU/adder/_239_ ) );
XNOR2_X1 \EXU/ALU/adder/_529_ ( .A(fanout_net_16 ), .B(\EXU/ALU/adder/_043_ ), .ZN(\EXU/ALU/adder/_240_ ) );
XNOR2_X1 \EXU/ALU/adder/_530_ ( .A(\EXU/ALU/adder/_240_ ), .B(\EXU/ALU/adder/_011_ ), .ZN(\EXU/ALU/adder/_241_ ) );
OR3_X1 \EXU/ALU/adder/_531_ ( .A1(\EXU/ALU/adder/_236_ ), .A2(\EXU/ALU/adder/_239_ ), .A3(\EXU/ALU/adder/_241_ ), .ZN(\EXU/ALU/adder/_242_ ) );
OAI21_X1 \EXU/ALU/adder/_532_ ( .A(\EXU/ALU/adder/_241_ ), .B1(\EXU/ALU/adder/_236_ ), .B2(\EXU/ALU/adder/_239_ ), .ZN(\EXU/ALU/adder/_243_ ) );
AND2_X1 \EXU/ALU/adder/_533_ ( .A1(\EXU/ALU/adder/_242_ ), .A2(\EXU/ALU/adder/_243_ ), .ZN(\EXU/ALU/adder/_076_ ) );
INV_X1 \EXU/ALU/adder/_534_ ( .A(\EXU/ALU/adder/_011_ ), .ZN(\EXU/ALU/adder/_244_ ) );
OR2_X1 \EXU/ALU/adder/_535_ ( .A1(\EXU/ALU/adder/_240_ ), .A2(\EXU/ALU/adder/_244_ ), .ZN(\EXU/ALU/adder/_245_ ) );
NAND2_X1 \EXU/ALU/adder/_536_ ( .A1(\EXU/ALU/adder/_243_ ), .A2(\EXU/ALU/adder/_245_ ), .ZN(\EXU/ALU/adder/_246_ ) );
XNOR2_X1 \EXU/ALU/adder/_537_ ( .A(fanout_net_16 ), .B(\EXU/ALU/adder/_044_ ), .ZN(\EXU/ALU/adder/_247_ ) );
XNOR2_X1 \EXU/ALU/adder/_538_ ( .A(\EXU/ALU/adder/_247_ ), .B(\EXU/ALU/adder/_012_ ), .ZN(\EXU/ALU/adder/_248_ ) );
INV_X1 \EXU/ALU/adder/_539_ ( .A(\EXU/ALU/adder/_248_ ), .ZN(\EXU/ALU/adder/_249_ ) );
XNOR2_X1 \EXU/ALU/adder/_540_ ( .A(\EXU/ALU/adder/_246_ ), .B(\EXU/ALU/adder/_249_ ), .ZN(\EXU/ALU/adder/_077_ ) );
AND2_X1 \EXU/ALU/adder/_541_ ( .A1(\EXU/ALU/adder/_241_ ), .A2(\EXU/ALU/adder/_248_ ), .ZN(\EXU/ALU/adder/_250_ ) );
AND2_X1 \EXU/ALU/adder/_542_ ( .A1(\EXU/ALU/adder/_234_ ), .A2(\EXU/ALU/adder/_250_ ), .ZN(\EXU/ALU/adder/_251_ ) );
INV_X1 \EXU/ALU/adder/_543_ ( .A(\EXU/ALU/adder/_251_ ), .ZN(\EXU/ALU/adder/_252_ ) );
OR2_X1 \EXU/ALU/adder/_544_ ( .A1(\EXU/ALU/adder/_224_ ), .A2(\EXU/ALU/adder/_252_ ), .ZN(\EXU/ALU/adder/_253_ ) );
OR2_X1 \EXU/ALU/adder/_545_ ( .A1(\EXU/ALU/adder/_249_ ), .A2(\EXU/ALU/adder/_245_ ), .ZN(\EXU/ALU/adder/_254_ ) );
INV_X1 \EXU/ALU/adder/_546_ ( .A(\EXU/ALU/adder/_012_ ), .ZN(\EXU/ALU/adder/_255_ ) );
OAI21_X1 \EXU/ALU/adder/_547_ ( .A(\EXU/ALU/adder/_254_ ), .B1(\EXU/ALU/adder/_255_ ), .B2(\EXU/ALU/adder/_247_ ), .ZN(\EXU/ALU/adder/_256_ ) );
AOI21_X1 \EXU/ALU/adder/_548_ ( .A(\EXU/ALU/adder/_256_ ), .B1(\EXU/ALU/adder/_239_ ), .B2(\EXU/ALU/adder/_250_ ), .ZN(\EXU/ALU/adder/_257_ ) );
AND2_X1 \EXU/ALU/adder/_549_ ( .A1(\EXU/ALU/adder/_253_ ), .A2(\EXU/ALU/adder/_257_ ), .ZN(\EXU/ALU/adder/_258_ ) );
XNOR2_X1 \EXU/ALU/adder/_550_ ( .A(fanout_net_16 ), .B(\EXU/ALU/adder/_046_ ), .ZN(\EXU/ALU/adder/_259_ ) );
XNOR2_X1 \EXU/ALU/adder/_551_ ( .A(\EXU/ALU/adder/_259_ ), .B(\EXU/ALU/adder/_014_ ), .ZN(\EXU/ALU/adder/_260_ ) );
XNOR2_X1 \EXU/ALU/adder/_552_ ( .A(\EXU/ALU/adder/_258_ ), .B(\EXU/ALU/adder/_260_ ), .ZN(\EXU/ALU/adder/_079_ ) );
INV_X1 \EXU/ALU/adder/_553_ ( .A(\EXU/ALU/adder/_260_ ), .ZN(\EXU/ALU/adder/_261_ ) );
OR2_X1 \EXU/ALU/adder/_554_ ( .A1(\EXU/ALU/adder/_258_ ), .A2(\EXU/ALU/adder/_261_ ), .ZN(\EXU/ALU/adder/_262_ ) );
INV_X1 \EXU/ALU/adder/_555_ ( .A(\EXU/ALU/adder/_014_ ), .ZN(\EXU/ALU/adder/_263_ ) );
OR2_X1 \EXU/ALU/adder/_556_ ( .A1(\EXU/ALU/adder/_259_ ), .A2(\EXU/ALU/adder/_263_ ), .ZN(\EXU/ALU/adder/_264_ ) );
NAND2_X1 \EXU/ALU/adder/_557_ ( .A1(\EXU/ALU/adder/_262_ ), .A2(\EXU/ALU/adder/_264_ ), .ZN(\EXU/ALU/adder/_265_ ) );
XNOR2_X1 \EXU/ALU/adder/_558_ ( .A(fanout_net_16 ), .B(\EXU/ALU/adder/_047_ ), .ZN(\EXU/ALU/adder/_266_ ) );
XNOR2_X1 \EXU/ALU/adder/_559_ ( .A(\EXU/ALU/adder/_266_ ), .B(\EXU/ALU/adder/_015_ ), .ZN(\EXU/ALU/adder/_267_ ) );
INV_X1 \EXU/ALU/adder/_560_ ( .A(\EXU/ALU/adder/_267_ ), .ZN(\EXU/ALU/adder/_268_ ) );
XNOR2_X1 \EXU/ALU/adder/_561_ ( .A(\EXU/ALU/adder/_265_ ), .B(\EXU/ALU/adder/_268_ ), .ZN(\EXU/ALU/adder/_080_ ) );
AOI211_X4 \EXU/ALU/adder/_562_ ( .A(\EXU/ALU/adder/_261_ ), .B(\EXU/ALU/adder/_268_ ), .C1(\EXU/ALU/adder/_253_ ), .C2(\EXU/ALU/adder/_257_ ), .ZN(\EXU/ALU/adder/_269_ ) );
OR2_X1 \EXU/ALU/adder/_563_ ( .A1(\EXU/ALU/adder/_268_ ), .A2(\EXU/ALU/adder/_264_ ), .ZN(\EXU/ALU/adder/_270_ ) );
INV_X1 \EXU/ALU/adder/_564_ ( .A(\EXU/ALU/adder/_015_ ), .ZN(\EXU/ALU/adder/_271_ ) );
OAI21_X1 \EXU/ALU/adder/_565_ ( .A(\EXU/ALU/adder/_270_ ), .B1(\EXU/ALU/adder/_271_ ), .B2(\EXU/ALU/adder/_266_ ), .ZN(\EXU/ALU/adder/_272_ ) );
NOR2_X1 \EXU/ALU/adder/_566_ ( .A1(\EXU/ALU/adder/_269_ ), .A2(\EXU/ALU/adder/_272_ ), .ZN(\EXU/ALU/adder/_273_ ) );
XNOR2_X1 \EXU/ALU/adder/_567_ ( .A(fanout_net_16 ), .B(\EXU/ALU/adder/_048_ ), .ZN(\EXU/ALU/adder/_274_ ) );
INV_X1 \EXU/ALU/adder/_568_ ( .A(\EXU/ALU/adder/_016_ ), .ZN(\EXU/ALU/adder/_275_ ) );
XNOR2_X1 \EXU/ALU/adder/_569_ ( .A(\EXU/ALU/adder/_274_ ), .B(\EXU/ALU/adder/_275_ ), .ZN(\EXU/ALU/adder/_276_ ) );
XOR2_X1 \EXU/ALU/adder/_570_ ( .A(\EXU/ALU/adder/_273_ ), .B(\EXU/ALU/adder/_276_ ), .Z(\EXU/ALU/adder/_081_ ) );
NOR2_X1 \EXU/ALU/adder/_571_ ( .A1(\EXU/ALU/adder/_273_ ), .A2(\EXU/ALU/adder/_276_ ), .ZN(\EXU/ALU/adder/_277_ ) );
NOR2_X1 \EXU/ALU/adder/_572_ ( .A1(\EXU/ALU/adder/_274_ ), .A2(\EXU/ALU/adder/_275_ ), .ZN(\EXU/ALU/adder/_278_ ) );
OR2_X1 \EXU/ALU/adder/_573_ ( .A1(\EXU/ALU/adder/_277_ ), .A2(\EXU/ALU/adder/_278_ ), .ZN(\EXU/ALU/adder/_279_ ) );
XNOR2_X1 \EXU/ALU/adder/_574_ ( .A(fanout_net_16 ), .B(\EXU/ALU/adder/_049_ ), .ZN(\EXU/ALU/adder/_280_ ) );
XNOR2_X1 \EXU/ALU/adder/_575_ ( .A(\EXU/ALU/adder/_280_ ), .B(\EXU/ALU/adder/_017_ ), .ZN(\EXU/ALU/adder/_281_ ) );
XNOR2_X1 \EXU/ALU/adder/_576_ ( .A(\EXU/ALU/adder/_279_ ), .B(\EXU/ALU/adder/_281_ ), .ZN(\EXU/ALU/adder/_282_ ) );
INV_X1 \EXU/ALU/adder/_577_ ( .A(\EXU/ALU/adder/_282_ ), .ZN(\EXU/ALU/adder/_082_ ) );
INV_X1 \EXU/ALU/adder/_578_ ( .A(\EXU/ALU/adder/_017_ ), .ZN(\EXU/ALU/adder/_283_ ) );
NOR2_X1 \EXU/ALU/adder/_579_ ( .A1(\EXU/ALU/adder/_280_ ), .A2(\EXU/ALU/adder/_283_ ), .ZN(\EXU/ALU/adder/_284_ ) );
AND2_X1 \EXU/ALU/adder/_580_ ( .A1(\EXU/ALU/adder/_280_ ), .A2(\EXU/ALU/adder/_283_ ), .ZN(\EXU/ALU/adder/_285_ ) );
NOR3_X1 \EXU/ALU/adder/_581_ ( .A1(\EXU/ALU/adder/_276_ ), .A2(\EXU/ALU/adder/_284_ ), .A3(\EXU/ALU/adder/_285_ ), .ZN(\EXU/ALU/adder/_286_ ) );
AND2_X1 \EXU/ALU/adder/_582_ ( .A1(\EXU/ALU/adder/_260_ ), .A2(\EXU/ALU/adder/_267_ ), .ZN(\EXU/ALU/adder/_287_ ) );
AND2_X1 \EXU/ALU/adder/_583_ ( .A1(\EXU/ALU/adder/_286_ ), .A2(\EXU/ALU/adder/_287_ ), .ZN(\EXU/ALU/adder/_288_ ) );
INV_X1 \EXU/ALU/adder/_584_ ( .A(\EXU/ALU/adder/_288_ ), .ZN(\EXU/ALU/adder/_289_ ) );
AOI211_X4 \EXU/ALU/adder/_585_ ( .A(\EXU/ALU/adder/_252_ ), .B(\EXU/ALU/adder/_289_ ), .C1(\EXU/ALU/adder/_217_ ), .C2(\EXU/ALU/adder/_223_ ), .ZN(\EXU/ALU/adder/_290_ ) );
NOR2_X1 \EXU/ALU/adder/_586_ ( .A1(\EXU/ALU/adder/_257_ ), .A2(\EXU/ALU/adder/_289_ ), .ZN(\EXU/ALU/adder/_291_ ) );
INV_X1 \EXU/ALU/adder/_587_ ( .A(\EXU/ALU/adder/_291_ ), .ZN(\EXU/ALU/adder/_292_ ) );
AOI221_X4 \EXU/ALU/adder/_588_ ( .A(\EXU/ALU/adder/_284_ ), .B1(\EXU/ALU/adder/_278_ ), .B2(\EXU/ALU/adder/_281_ ), .C1(\EXU/ALU/adder/_272_ ), .C2(\EXU/ALU/adder/_286_ ), .ZN(\EXU/ALU/adder/_293_ ) );
AND2_X1 \EXU/ALU/adder/_589_ ( .A1(\EXU/ALU/adder/_292_ ), .A2(\EXU/ALU/adder/_293_ ), .ZN(\EXU/ALU/adder/_294_ ) );
INV_X1 \EXU/ALU/adder/_590_ ( .A(\EXU/ALU/adder/_294_ ), .ZN(\EXU/ALU/adder/_295_ ) );
XNOR2_X1 \EXU/ALU/adder/_591_ ( .A(fanout_net_16 ), .B(\EXU/ALU/adder/_050_ ), .ZN(\EXU/ALU/adder/_296_ ) );
XNOR2_X1 \EXU/ALU/adder/_592_ ( .A(\EXU/ALU/adder/_296_ ), .B(\EXU/ALU/adder/_018_ ), .ZN(\EXU/ALU/adder/_297_ ) );
OR3_X1 \EXU/ALU/adder/_593_ ( .A1(\EXU/ALU/adder/_290_ ), .A2(\EXU/ALU/adder/_295_ ), .A3(\EXU/ALU/adder/_297_ ), .ZN(\EXU/ALU/adder/_298_ ) );
OAI21_X1 \EXU/ALU/adder/_594_ ( .A(\EXU/ALU/adder/_297_ ), .B1(\EXU/ALU/adder/_290_ ), .B2(\EXU/ALU/adder/_295_ ), .ZN(\EXU/ALU/adder/_299_ ) );
AND2_X1 \EXU/ALU/adder/_595_ ( .A1(\EXU/ALU/adder/_298_ ), .A2(\EXU/ALU/adder/_299_ ), .ZN(\EXU/ALU/adder/_083_ ) );
INV_X1 \EXU/ALU/adder/_596_ ( .A(\EXU/ALU/adder/_018_ ), .ZN(\EXU/ALU/adder/_300_ ) );
NOR2_X1 \EXU/ALU/adder/_597_ ( .A1(\EXU/ALU/adder/_296_ ), .A2(\EXU/ALU/adder/_300_ ), .ZN(\EXU/ALU/adder/_301_ ) );
INV_X1 \EXU/ALU/adder/_598_ ( .A(\EXU/ALU/adder/_301_ ), .ZN(\EXU/ALU/adder/_302_ ) );
AND2_X1 \EXU/ALU/adder/_599_ ( .A1(\EXU/ALU/adder/_299_ ), .A2(\EXU/ALU/adder/_302_ ), .ZN(\EXU/ALU/adder/_303_ ) );
XNOR2_X1 \EXU/ALU/adder/_600_ ( .A(fanout_net_16 ), .B(\EXU/ALU/adder/_051_ ), .ZN(\EXU/ALU/adder/_304_ ) );
XNOR2_X1 \EXU/ALU/adder/_601_ ( .A(\EXU/ALU/adder/_304_ ), .B(\EXU/ALU/adder/_019_ ), .ZN(\EXU/ALU/adder/_305_ ) );
XNOR2_X1 \EXU/ALU/adder/_602_ ( .A(\EXU/ALU/adder/_303_ ), .B(\EXU/ALU/adder/_305_ ), .ZN(\EXU/ALU/adder/_084_ ) );
AND2_X1 \EXU/ALU/adder/_603_ ( .A1(\EXU/ALU/adder/_297_ ), .A2(\EXU/ALU/adder/_305_ ), .ZN(\EXU/ALU/adder/_306_ ) );
OAI21_X1 \EXU/ALU/adder/_604_ ( .A(\EXU/ALU/adder/_306_ ), .B1(\EXU/ALU/adder/_290_ ), .B2(\EXU/ALU/adder/_295_ ), .ZN(\EXU/ALU/adder/_307_ ) );
NAND2_X1 \EXU/ALU/adder/_605_ ( .A1(\EXU/ALU/adder/_305_ ), .A2(\EXU/ALU/adder/_301_ ), .ZN(\EXU/ALU/adder/_308_ ) );
INV_X1 \EXU/ALU/adder/_606_ ( .A(\EXU/ALU/adder/_019_ ), .ZN(\EXU/ALU/adder/_309_ ) );
OAI21_X1 \EXU/ALU/adder/_607_ ( .A(\EXU/ALU/adder/_308_ ), .B1(\EXU/ALU/adder/_309_ ), .B2(\EXU/ALU/adder/_304_ ), .ZN(\EXU/ALU/adder/_310_ ) );
INV_X1 \EXU/ALU/adder/_608_ ( .A(\EXU/ALU/adder/_310_ ), .ZN(\EXU/ALU/adder/_311_ ) );
XNOR2_X1 \EXU/ALU/adder/_609_ ( .A(fanout_net_16 ), .B(\EXU/ALU/adder/_052_ ), .ZN(\EXU/ALU/adder/_312_ ) );
XNOR2_X1 \EXU/ALU/adder/_610_ ( .A(\EXU/ALU/adder/_312_ ), .B(\EXU/ALU/adder/_020_ ), .ZN(\EXU/ALU/adder/_313_ ) );
INV_X1 \EXU/ALU/adder/_611_ ( .A(\EXU/ALU/adder/_313_ ), .ZN(\EXU/ALU/adder/_314_ ) );
AND3_X1 \EXU/ALU/adder/_612_ ( .A1(\EXU/ALU/adder/_307_ ), .A2(\EXU/ALU/adder/_311_ ), .A3(\EXU/ALU/adder/_314_ ), .ZN(\EXU/ALU/adder/_315_ ) );
AOI21_X1 \EXU/ALU/adder/_613_ ( .A(\EXU/ALU/adder/_314_ ), .B1(\EXU/ALU/adder/_307_ ), .B2(\EXU/ALU/adder/_311_ ), .ZN(\EXU/ALU/adder/_316_ ) );
NOR2_X1 \EXU/ALU/adder/_614_ ( .A1(\EXU/ALU/adder/_315_ ), .A2(\EXU/ALU/adder/_316_ ), .ZN(\EXU/ALU/adder/_085_ ) );
INV_X1 \EXU/ALU/adder/_615_ ( .A(\EXU/ALU/adder/_020_ ), .ZN(\EXU/ALU/adder/_317_ ) );
NOR2_X1 \EXU/ALU/adder/_616_ ( .A1(\EXU/ALU/adder/_312_ ), .A2(\EXU/ALU/adder/_317_ ), .ZN(\EXU/ALU/adder/_318_ ) );
OR2_X1 \EXU/ALU/adder/_617_ ( .A1(\EXU/ALU/adder/_316_ ), .A2(\EXU/ALU/adder/_318_ ), .ZN(\EXU/ALU/adder/_319_ ) );
XNOR2_X1 \EXU/ALU/adder/_618_ ( .A(fanout_net_16 ), .B(\EXU/ALU/adder/_053_ ), .ZN(\EXU/ALU/adder/_320_ ) );
XNOR2_X1 \EXU/ALU/adder/_619_ ( .A(\EXU/ALU/adder/_320_ ), .B(\EXU/ALU/adder/_021_ ), .ZN(\EXU/ALU/adder/_321_ ) );
XNOR2_X1 \EXU/ALU/adder/_620_ ( .A(\EXU/ALU/adder/_319_ ), .B(\EXU/ALU/adder/_321_ ), .ZN(\EXU/ALU/adder/_322_ ) );
INV_X1 \EXU/ALU/adder/_621_ ( .A(\EXU/ALU/adder/_322_ ), .ZN(\EXU/ALU/adder/_086_ ) );
AND2_X1 \EXU/ALU/adder/_622_ ( .A1(\EXU/ALU/adder/_313_ ), .A2(\EXU/ALU/adder/_321_ ), .ZN(\EXU/ALU/adder/_323_ ) );
OAI211_X2 \EXU/ALU/adder/_623_ ( .A(\EXU/ALU/adder/_306_ ), .B(\EXU/ALU/adder/_323_ ), .C1(\EXU/ALU/adder/_290_ ), .C2(\EXU/ALU/adder/_295_ ), .ZN(\EXU/ALU/adder/_324_ ) );
NAND2_X1 \EXU/ALU/adder/_624_ ( .A1(\EXU/ALU/adder/_321_ ), .A2(\EXU/ALU/adder/_318_ ), .ZN(\EXU/ALU/adder/_325_ ) );
INV_X1 \EXU/ALU/adder/_625_ ( .A(\EXU/ALU/adder/_021_ ), .ZN(\EXU/ALU/adder/_326_ ) );
OAI21_X1 \EXU/ALU/adder/_626_ ( .A(\EXU/ALU/adder/_325_ ), .B1(\EXU/ALU/adder/_326_ ), .B2(\EXU/ALU/adder/_320_ ), .ZN(\EXU/ALU/adder/_327_ ) );
AOI21_X1 \EXU/ALU/adder/_627_ ( .A(\EXU/ALU/adder/_327_ ), .B1(\EXU/ALU/adder/_310_ ), .B2(\EXU/ALU/adder/_323_ ), .ZN(\EXU/ALU/adder/_328_ ) );
XNOR2_X1 \EXU/ALU/adder/_628_ ( .A(fanout_net_16 ), .B(\EXU/ALU/adder/_054_ ), .ZN(\EXU/ALU/adder/_329_ ) );
XNOR2_X1 \EXU/ALU/adder/_629_ ( .A(\EXU/ALU/adder/_329_ ), .B(\EXU/ALU/adder/_022_ ), .ZN(\EXU/ALU/adder/_330_ ) );
INV_X1 \EXU/ALU/adder/_630_ ( .A(\EXU/ALU/adder/_330_ ), .ZN(\EXU/ALU/adder/_331_ ) );
AND3_X1 \EXU/ALU/adder/_631_ ( .A1(\EXU/ALU/adder/_324_ ), .A2(\EXU/ALU/adder/_328_ ), .A3(\EXU/ALU/adder/_331_ ), .ZN(\EXU/ALU/adder/_332_ ) );
AOI21_X1 \EXU/ALU/adder/_632_ ( .A(\EXU/ALU/adder/_331_ ), .B1(\EXU/ALU/adder/_324_ ), .B2(\EXU/ALU/adder/_328_ ), .ZN(\EXU/ALU/adder/_333_ ) );
NOR2_X1 \EXU/ALU/adder/_633_ ( .A1(\EXU/ALU/adder/_332_ ), .A2(\EXU/ALU/adder/_333_ ), .ZN(\EXU/ALU/adder/_087_ ) );
INV_X1 \EXU/ALU/adder/_634_ ( .A(\EXU/ALU/adder/_022_ ), .ZN(\EXU/ALU/adder/_334_ ) );
NOR2_X1 \EXU/ALU/adder/_635_ ( .A1(\EXU/ALU/adder/_329_ ), .A2(\EXU/ALU/adder/_334_ ), .ZN(\EXU/ALU/adder/_335_ ) );
OR2_X1 \EXU/ALU/adder/_636_ ( .A1(\EXU/ALU/adder/_333_ ), .A2(\EXU/ALU/adder/_335_ ), .ZN(\EXU/ALU/adder/_336_ ) );
XNOR2_X1 \EXU/ALU/adder/_637_ ( .A(fanout_net_16 ), .B(\EXU/ALU/adder/_055_ ), .ZN(\EXU/ALU/adder/_337_ ) );
XNOR2_X1 \EXU/ALU/adder/_638_ ( .A(\EXU/ALU/adder/_337_ ), .B(\EXU/ALU/adder/_023_ ), .ZN(\EXU/ALU/adder/_338_ ) );
XNOR2_X1 \EXU/ALU/adder/_639_ ( .A(\EXU/ALU/adder/_336_ ), .B(\EXU/ALU/adder/_338_ ), .ZN(\EXU/ALU/adder/_339_ ) );
INV_X1 \EXU/ALU/adder/_640_ ( .A(\EXU/ALU/adder/_339_ ), .ZN(\EXU/ALU/adder/_088_ ) );
AND2_X1 \EXU/ALU/adder/_641_ ( .A1(\EXU/ALU/adder/_333_ ), .A2(\EXU/ALU/adder/_338_ ), .ZN(\EXU/ALU/adder/_340_ ) );
NAND2_X1 \EXU/ALU/adder/_642_ ( .A1(\EXU/ALU/adder/_338_ ), .A2(\EXU/ALU/adder/_335_ ), .ZN(\EXU/ALU/adder/_341_ ) );
INV_X1 \EXU/ALU/adder/_643_ ( .A(\EXU/ALU/adder/_023_ ), .ZN(\EXU/ALU/adder/_342_ ) );
OAI21_X1 \EXU/ALU/adder/_644_ ( .A(\EXU/ALU/adder/_341_ ), .B1(\EXU/ALU/adder/_342_ ), .B2(\EXU/ALU/adder/_337_ ), .ZN(\EXU/ALU/adder/_343_ ) );
XNOR2_X1 \EXU/ALU/adder/_645_ ( .A(\EXU/ALU/adder/_000_ ), .B(\EXU/ALU/adder/_057_ ), .ZN(\EXU/ALU/adder/_344_ ) );
XNOR2_X1 \EXU/ALU/adder/_646_ ( .A(\EXU/ALU/adder/_344_ ), .B(\EXU/ALU/adder/_025_ ), .ZN(\EXU/ALU/adder/_345_ ) );
OR3_X1 \EXU/ALU/adder/_647_ ( .A1(\EXU/ALU/adder/_340_ ), .A2(\EXU/ALU/adder/_343_ ), .A3(\EXU/ALU/adder/_345_ ), .ZN(\EXU/ALU/adder/_346_ ) );
OAI21_X1 \EXU/ALU/adder/_648_ ( .A(\EXU/ALU/adder/_345_ ), .B1(\EXU/ALU/adder/_340_ ), .B2(\EXU/ALU/adder/_343_ ), .ZN(\EXU/ALU/adder/_347_ ) );
AND2_X1 \EXU/ALU/adder/_649_ ( .A1(\EXU/ALU/adder/_346_ ), .A2(\EXU/ALU/adder/_347_ ), .ZN(\EXU/ALU/adder/_090_ ) );
INV_X1 \EXU/ALU/adder/_650_ ( .A(\EXU/ALU/adder/_025_ ), .ZN(\EXU/ALU/adder/_348_ ) );
NOR2_X1 \EXU/ALU/adder/_651_ ( .A1(\EXU/ALU/adder/_344_ ), .A2(\EXU/ALU/adder/_348_ ), .ZN(\EXU/ALU/adder/_349_ ) );
INV_X1 \EXU/ALU/adder/_652_ ( .A(\EXU/ALU/adder/_349_ ), .ZN(\EXU/ALU/adder/_350_ ) );
NAND2_X1 \EXU/ALU/adder/_653_ ( .A1(\EXU/ALU/adder/_347_ ), .A2(\EXU/ALU/adder/_350_ ), .ZN(\EXU/ALU/adder/_351_ ) );
XNOR2_X1 \EXU/ALU/adder/_654_ ( .A(\EXU/ALU/adder/_000_ ), .B(\EXU/ALU/adder/_058_ ), .ZN(\EXU/ALU/adder/_352_ ) );
XNOR2_X1 \EXU/ALU/adder/_655_ ( .A(\EXU/ALU/adder/_352_ ), .B(\EXU/ALU/adder/_026_ ), .ZN(\EXU/ALU/adder/_353_ ) );
XOR2_X1 \EXU/ALU/adder/_656_ ( .A(\EXU/ALU/adder/_351_ ), .B(\EXU/ALU/adder/_353_ ), .Z(\EXU/ALU/adder/_091_ ) );
OR4_X4 \EXU/ALU/adder/_657_ ( .A1(\EXU/ALU/adder/_098_ ), .A2(\EXU/ALU/adder/_074_ ), .A3(\EXU/ALU/adder/_070_ ), .A4(\EXU/ALU/adder/_068_ ), .ZN(\EXU/ALU/adder/_354_ ) );
OR3_X2 \EXU/ALU/adder/_658_ ( .A1(\EXU/ALU/adder/_089_ ), .A2(\EXU/ALU/adder/_067_ ), .A3(\EXU/ALU/adder/_078_ ), .ZN(\EXU/ALU/adder/_355_ ) );
OR3_X1 \EXU/ALU/adder/_659_ ( .A1(\EXU/ALU/adder/_093_ ), .A2(\EXU/ALU/adder/_092_ ), .A3(\EXU/ALU/adder/_355_ ), .ZN(\EXU/ALU/adder/_356_ ) );
OR4_X4 \EXU/ALU/adder/_660_ ( .A1(\EXU/ALU/adder/_094_ ), .A2(\EXU/ALU/adder/_095_ ), .A3(\EXU/ALU/adder/_097_ ), .A4(\EXU/ALU/adder/_356_ ), .ZN(\EXU/ALU/adder/_357_ ) );
OR3_X4 \EXU/ALU/adder/_661_ ( .A1(\EXU/ALU/adder/_354_ ), .A2(\EXU/ALU/adder/_096_ ), .A3(\EXU/ALU/adder/_357_ ), .ZN(\EXU/ALU/adder/_358_ ) );
OR3_X4 \EXU/ALU/adder/_662_ ( .A1(\EXU/ALU/adder/_358_ ), .A2(\EXU/ALU/adder/_069_ ), .A3(\EXU/ALU/adder/_072_ ), .ZN(\EXU/ALU/adder/_359_ ) );
NOR3_X4 \EXU/ALU/adder/_663_ ( .A1(\EXU/ALU/adder/_359_ ), .A2(\EXU/ALU/adder/_071_ ), .A3(\EXU/ALU/adder/_075_ ), .ZN(\EXU/ALU/adder/_360_ ) );
NOR4_X1 \EXU/ALU/adder/_664_ ( .A1(\EXU/ALU/adder/_080_ ), .A2(\EXU/ALU/adder/_076_ ), .A3(\EXU/ALU/adder/_079_ ), .A4(\EXU/ALU/adder/_083_ ), .ZN(\EXU/ALU/adder/_361_ ) );
NAND2_X1 \EXU/ALU/adder/_665_ ( .A1(\EXU/ALU/adder/_360_ ), .A2(\EXU/ALU/adder/_361_ ), .ZN(\EXU/ALU/adder/_362_ ) );
OR2_X1 \EXU/ALU/adder/_666_ ( .A1(\EXU/ALU/adder/_081_ ), .A2(\EXU/ALU/adder/_085_ ), .ZN(\EXU/ALU/adder/_363_ ) );
OR4_X2 \EXU/ALU/adder/_667_ ( .A1(\EXU/ALU/adder/_084_ ), .A2(\EXU/ALU/adder/_362_ ), .A3(\EXU/ALU/adder/_087_ ), .A4(\EXU/ALU/adder/_363_ ), .ZN(\EXU/ALU/adder/_364_ ) );
OR3_X4 \EXU/ALU/adder/_668_ ( .A1(\EXU/ALU/adder/_364_ ), .A2(\EXU/ALU/adder/_086_ ), .A3(\EXU/ALU/adder/_090_ ), .ZN(\EXU/ALU/adder/_365_ ) );
OR4_X4 \EXU/ALU/adder/_669_ ( .A1(\EXU/ALU/adder/_073_ ), .A2(\EXU/ALU/adder/_365_ ), .A3(\EXU/ALU/adder/_077_ ), .A4(\EXU/ALU/adder/_082_ ), .ZN(\EXU/ALU/adder/_366_ ) );
NOR3_X1 \EXU/ALU/adder/_670_ ( .A1(\EXU/ALU/adder/_366_ ), .A2(\EXU/ALU/adder/_088_ ), .A3(\EXU/ALU/adder/_091_ ), .ZN(\EXU/ALU/adder/_099_ ) );
XNOR2_X1 \EXU/ALU/adder/_671_ ( .A(\EXU/ALU/adder/_091_ ), .B(\EXU/ALU/adder/_026_ ), .ZN(\EXU/ALU/adder/_367_ ) );
NOR2_X1 \EXU/ALU/adder/_672_ ( .A1(\EXU/ALU/adder/_367_ ), .A2(\EXU/ALU/adder/_353_ ), .ZN(\EXU/ALU/adder/_066_ ) );
OAI211_X2 \EXU/ALU/adder/_673_ ( .A(\EXU/ALU/adder/_345_ ), .B(\EXU/ALU/adder/_353_ ), .C1(\EXU/ALU/adder/_340_ ), .C2(\EXU/ALU/adder/_343_ ), .ZN(\EXU/ALU/adder/_368_ ) );
NAND2_X1 \EXU/ALU/adder/_674_ ( .A1(\EXU/ALU/adder/_353_ ), .A2(\EXU/ALU/adder/_349_ ), .ZN(\EXU/ALU/adder/_369_ ) );
INV_X1 \EXU/ALU/adder/_675_ ( .A(\EXU/ALU/adder/_026_ ), .ZN(\EXU/ALU/adder/_370_ ) );
OAI211_X2 \EXU/ALU/adder/_676_ ( .A(\EXU/ALU/adder/_368_ ), .B(\EXU/ALU/adder/_369_ ), .C1(\EXU/ALU/adder/_370_ ), .C2(\EXU/ALU/adder/_352_ ), .ZN(\EXU/ALU/adder/_001_ ) );
BUF_X1 \EXU/ALU/adder/_677_ ( .A(\EXU/casez_tmp_0 [0] ), .Z(\EXU/ALU/adder/_034_ ) );
BUF_X1 \EXU/ALU/adder/_678_ ( .A(\EXU/ALU/_aluControl_io_isSub ), .Z(\EXU/ALU/adder/_000_ ) );
BUF_X1 \EXU/ALU/adder/_679_ ( .A(\EXU/_0000_ ), .Z(\EXU/ALU/adder/_002_ ) );
BUF_X1 \EXU/ALU/adder/_680_ ( .A(\EXU/ALU/adder/_067_ ), .Z(\EXU/ALU/_adder_io_result [0] ) );
BUF_X1 \EXU/ALU/adder/_681_ ( .A(\EXU/casez_tmp_0 [1] ), .Z(\EXU/ALU/adder/_045_ ) );
BUF_X1 \EXU/ALU/adder/_682_ ( .A(\EXU/_0011_ ), .Z(\EXU/ALU/adder/_013_ ) );
BUF_X1 \EXU/ALU/adder/_683_ ( .A(\EXU/ALU/adder/_078_ ), .Z(\EXU/ALU/_adder_io_result [1] ) );
BUF_X1 \EXU/ALU/adder/_684_ ( .A(\EXU/casez_tmp_0 [2] ), .Z(\EXU/ALU/adder/_056_ ) );
BUF_X1 \EXU/ALU/adder/_685_ ( .A(\EXU/_0022_ ), .Z(\EXU/ALU/adder/_024_ ) );
BUF_X1 \EXU/ALU/adder/_686_ ( .A(\EXU/ALU/adder/_089_ ), .Z(\EXU/ALU/_adder_io_result [2] ) );
BUF_X1 \EXU/ALU/adder/_687_ ( .A(\EXU/casez_tmp_0 [3] ), .Z(\EXU/ALU/adder/_059_ ) );
BUF_X1 \EXU/ALU/adder/_688_ ( .A(\EXU/_0025_ ), .Z(\EXU/ALU/adder/_027_ ) );
BUF_X1 \EXU/ALU/adder/_689_ ( .A(\EXU/ALU/adder/_092_ ), .Z(\EXU/ALU/_adder_io_result [3] ) );
BUF_X1 \EXU/ALU/adder/_690_ ( .A(\EXU/casez_tmp_0 [4] ), .Z(\EXU/ALU/adder/_060_ ) );
BUF_X1 \EXU/ALU/adder/_691_ ( .A(\EXU/_0026_ ), .Z(\EXU/ALU/adder/_028_ ) );
BUF_X1 \EXU/ALU/adder/_692_ ( .A(\EXU/ALU/adder/_093_ ), .Z(\EXU/ALU/_adder_io_result [4] ) );
BUF_X1 \EXU/ALU/adder/_693_ ( .A(\EXU/casez_tmp_0 [5] ), .Z(\EXU/ALU/adder/_061_ ) );
BUF_X1 \EXU/ALU/adder/_694_ ( .A(\EXU/_0027_ ), .Z(\EXU/ALU/adder/_029_ ) );
BUF_X1 \EXU/ALU/adder/_695_ ( .A(\EXU/ALU/adder/_094_ ), .Z(\EXU/ALU/_adder_io_result [5] ) );
BUF_X1 \EXU/ALU/adder/_696_ ( .A(\EXU/casez_tmp_0 [6] ), .Z(\EXU/ALU/adder/_062_ ) );
BUF_X1 \EXU/ALU/adder/_697_ ( .A(\EXU/_0028_ ), .Z(\EXU/ALU/adder/_030_ ) );
BUF_X1 \EXU/ALU/adder/_698_ ( .A(\EXU/ALU/adder/_095_ ), .Z(\EXU/ALU/_adder_io_result [6] ) );
BUF_X1 \EXU/ALU/adder/_699_ ( .A(\EXU/casez_tmp_0 [7] ), .Z(\EXU/ALU/adder/_063_ ) );
BUF_X1 \EXU/ALU/adder/_700_ ( .A(\EXU/_0029_ ), .Z(\EXU/ALU/adder/_031_ ) );
BUF_X1 \EXU/ALU/adder/_701_ ( .A(\EXU/ALU/adder/_096_ ), .Z(\EXU/ALU/_adder_io_result [7] ) );
BUF_X1 \EXU/ALU/adder/_702_ ( .A(\EXU/casez_tmp_0 [8] ), .Z(\EXU/ALU/adder/_064_ ) );
BUF_X1 \EXU/ALU/adder/_703_ ( .A(\EXU/_0030_ ), .Z(\EXU/ALU/adder/_032_ ) );
BUF_X1 \EXU/ALU/adder/_704_ ( .A(\EXU/ALU/adder/_097_ ), .Z(\EXU/ALU/_adder_io_result [8] ) );
BUF_X1 \EXU/ALU/adder/_705_ ( .A(\EXU/casez_tmp_0 [9] ), .Z(\EXU/ALU/adder/_065_ ) );
BUF_X1 \EXU/ALU/adder/_706_ ( .A(\EXU/_0031_ ), .Z(\EXU/ALU/adder/_033_ ) );
BUF_X1 \EXU/ALU/adder/_707_ ( .A(\EXU/ALU/adder/_098_ ), .Z(\EXU/ALU/_adder_io_result [9] ) );
BUF_X1 \EXU/ALU/adder/_708_ ( .A(\EXU/casez_tmp_0 [10] ), .Z(\EXU/ALU/adder/_035_ ) );
BUF_X1 \EXU/ALU/adder/_709_ ( .A(\EXU/_0001_ ), .Z(\EXU/ALU/adder/_003_ ) );
BUF_X1 \EXU/ALU/adder/_710_ ( .A(\EXU/ALU/adder/_068_ ), .Z(\EXU/ALU/_adder_io_result [10] ) );
BUF_X1 \EXU/ALU/adder/_711_ ( .A(\EXU/casez_tmp_0 [11] ), .Z(\EXU/ALU/adder/_036_ ) );
BUF_X1 \EXU/ALU/adder/_712_ ( .A(\EXU/_0002_ ), .Z(\EXU/ALU/adder/_004_ ) );
BUF_X1 \EXU/ALU/adder/_713_ ( .A(\EXU/ALU/adder/_069_ ), .Z(\EXU/ALU/_adder_io_result [11] ) );
BUF_X1 \EXU/ALU/adder/_714_ ( .A(\EXU/casez_tmp_0 [12] ), .Z(\EXU/ALU/adder/_037_ ) );
BUF_X1 \EXU/ALU/adder/_715_ ( .A(\EXU/_0003_ ), .Z(\EXU/ALU/adder/_005_ ) );
BUF_X1 \EXU/ALU/adder/_716_ ( .A(\EXU/ALU/adder/_070_ ), .Z(\EXU/ALU/_adder_io_result [12] ) );
BUF_X1 \EXU/ALU/adder/_717_ ( .A(\EXU/casez_tmp_0 [13] ), .Z(\EXU/ALU/adder/_038_ ) );
BUF_X1 \EXU/ALU/adder/_718_ ( .A(\EXU/_0004_ ), .Z(\EXU/ALU/adder/_006_ ) );
BUF_X1 \EXU/ALU/adder/_719_ ( .A(\EXU/ALU/adder/_071_ ), .Z(\EXU/ALU/_adder_io_result [13] ) );
BUF_X1 \EXU/ALU/adder/_720_ ( .A(\EXU/casez_tmp_0 [14] ), .Z(\EXU/ALU/adder/_039_ ) );
BUF_X1 \EXU/ALU/adder/_721_ ( .A(\EXU/_0005_ ), .Z(\EXU/ALU/adder/_007_ ) );
BUF_X1 \EXU/ALU/adder/_722_ ( .A(\EXU/ALU/adder/_072_ ), .Z(\EXU/ALU/_adder_io_result [14] ) );
BUF_X1 \EXU/ALU/adder/_723_ ( .A(\EXU/casez_tmp_0 [15] ), .Z(\EXU/ALU/adder/_040_ ) );
BUF_X1 \EXU/ALU/adder/_724_ ( .A(\EXU/_0006_ ), .Z(\EXU/ALU/adder/_008_ ) );
BUF_X1 \EXU/ALU/adder/_725_ ( .A(\EXU/ALU/adder/_073_ ), .Z(\EXU/ALU/_adder_io_result [15] ) );
BUF_X1 \EXU/ALU/adder/_726_ ( .A(\EXU/casez_tmp_0 [16] ), .Z(\EXU/ALU/adder/_041_ ) );
BUF_X1 \EXU/ALU/adder/_727_ ( .A(\EXU/_0007_ ), .Z(\EXU/ALU/adder/_009_ ) );
BUF_X1 \EXU/ALU/adder/_728_ ( .A(\EXU/ALU/adder/_074_ ), .Z(\EXU/ALU/_adder_io_result [16] ) );
BUF_X1 \EXU/ALU/adder/_729_ ( .A(\EXU/_0008_ ), .Z(\EXU/ALU/adder/_010_ ) );
BUF_X1 \EXU/ALU/adder/_730_ ( .A(\EXU/casez_tmp_0 [17] ), .Z(\EXU/ALU/adder/_042_ ) );
BUF_X1 \EXU/ALU/adder/_731_ ( .A(\EXU/ALU/adder/_075_ ), .Z(\EXU/ALU/_adder_io_result [17] ) );
BUF_X1 \EXU/ALU/adder/_732_ ( .A(\EXU/casez_tmp_0 [18] ), .Z(\EXU/ALU/adder/_043_ ) );
BUF_X1 \EXU/ALU/adder/_733_ ( .A(\EXU/_0009_ ), .Z(\EXU/ALU/adder/_011_ ) );
BUF_X1 \EXU/ALU/adder/_734_ ( .A(\EXU/ALU/adder/_076_ ), .Z(\EXU/ALU/_adder_io_result [18] ) );
BUF_X1 \EXU/ALU/adder/_735_ ( .A(\EXU/casez_tmp_0 [19] ), .Z(\EXU/ALU/adder/_044_ ) );
BUF_X1 \EXU/ALU/adder/_736_ ( .A(\EXU/_0010_ ), .Z(\EXU/ALU/adder/_012_ ) );
BUF_X1 \EXU/ALU/adder/_737_ ( .A(\EXU/ALU/adder/_077_ ), .Z(\EXU/ALU/_adder_io_result [19] ) );
BUF_X1 \EXU/ALU/adder/_738_ ( .A(\EXU/casez_tmp_0 [20] ), .Z(\EXU/ALU/adder/_046_ ) );
BUF_X1 \EXU/ALU/adder/_739_ ( .A(\EXU/_0012_ ), .Z(\EXU/ALU/adder/_014_ ) );
BUF_X1 \EXU/ALU/adder/_740_ ( .A(\EXU/ALU/adder/_079_ ), .Z(\EXU/ALU/_adder_io_result [20] ) );
BUF_X1 \EXU/ALU/adder/_741_ ( .A(\EXU/_0013_ ), .Z(\EXU/ALU/adder/_015_ ) );
BUF_X1 \EXU/ALU/adder/_742_ ( .A(\EXU/casez_tmp_0 [21] ), .Z(\EXU/ALU/adder/_047_ ) );
BUF_X1 \EXU/ALU/adder/_743_ ( .A(\EXU/ALU/adder/_080_ ), .Z(\EXU/ALU/_adder_io_result [21] ) );
BUF_X1 \EXU/ALU/adder/_744_ ( .A(\EXU/casez_tmp_0 [22] ), .Z(\EXU/ALU/adder/_048_ ) );
BUF_X1 \EXU/ALU/adder/_745_ ( .A(\EXU/_0014_ ), .Z(\EXU/ALU/adder/_016_ ) );
BUF_X1 \EXU/ALU/adder/_746_ ( .A(\EXU/ALU/adder/_081_ ), .Z(\EXU/ALU/_adder_io_result [22] ) );
BUF_X1 \EXU/ALU/adder/_747_ ( .A(\EXU/casez_tmp_0 [23] ), .Z(\EXU/ALU/adder/_049_ ) );
BUF_X1 \EXU/ALU/adder/_748_ ( .A(\EXU/_0015_ ), .Z(\EXU/ALU/adder/_017_ ) );
BUF_X1 \EXU/ALU/adder/_749_ ( .A(\EXU/ALU/adder/_082_ ), .Z(\EXU/ALU/_adder_io_result [23] ) );
BUF_X1 \EXU/ALU/adder/_750_ ( .A(\EXU/casez_tmp_0 [24] ), .Z(\EXU/ALU/adder/_050_ ) );
BUF_X1 \EXU/ALU/adder/_751_ ( .A(\EXU/_0016_ ), .Z(\EXU/ALU/adder/_018_ ) );
BUF_X1 \EXU/ALU/adder/_752_ ( .A(\EXU/ALU/adder/_083_ ), .Z(\EXU/ALU/_adder_io_result [24] ) );
BUF_X1 \EXU/ALU/adder/_753_ ( .A(\EXU/casez_tmp_0 [25] ), .Z(\EXU/ALU/adder/_051_ ) );
BUF_X1 \EXU/ALU/adder/_754_ ( .A(\EXU/_0017_ ), .Z(\EXU/ALU/adder/_019_ ) );
BUF_X1 \EXU/ALU/adder/_755_ ( .A(\EXU/ALU/adder/_084_ ), .Z(\EXU/ALU/_adder_io_result [25] ) );
BUF_X1 \EXU/ALU/adder/_756_ ( .A(\EXU/casez_tmp_0 [26] ), .Z(\EXU/ALU/adder/_052_ ) );
BUF_X1 \EXU/ALU/adder/_757_ ( .A(\EXU/_0018_ ), .Z(\EXU/ALU/adder/_020_ ) );
BUF_X1 \EXU/ALU/adder/_758_ ( .A(\EXU/ALU/adder/_085_ ), .Z(\EXU/ALU/_adder_io_result [26] ) );
BUF_X1 \EXU/ALU/adder/_759_ ( .A(\EXU/casez_tmp_0 [27] ), .Z(\EXU/ALU/adder/_053_ ) );
BUF_X1 \EXU/ALU/adder/_760_ ( .A(\EXU/_0019_ ), .Z(\EXU/ALU/adder/_021_ ) );
BUF_X1 \EXU/ALU/adder/_761_ ( .A(\EXU/ALU/adder/_086_ ), .Z(\EXU/ALU/_adder_io_result [27] ) );
BUF_X1 \EXU/ALU/adder/_762_ ( .A(\EXU/casez_tmp_0 [28] ), .Z(\EXU/ALU/adder/_054_ ) );
BUF_X1 \EXU/ALU/adder/_763_ ( .A(\EXU/_0020_ ), .Z(\EXU/ALU/adder/_022_ ) );
BUF_X1 \EXU/ALU/adder/_764_ ( .A(\EXU/ALU/adder/_087_ ), .Z(\EXU/ALU/_adder_io_result [28] ) );
BUF_X1 \EXU/ALU/adder/_765_ ( .A(\EXU/casez_tmp_0 [29] ), .Z(\EXU/ALU/adder/_055_ ) );
BUF_X1 \EXU/ALU/adder/_766_ ( .A(\EXU/_0021_ ), .Z(\EXU/ALU/adder/_023_ ) );
BUF_X1 \EXU/ALU/adder/_767_ ( .A(\EXU/ALU/adder/_088_ ), .Z(\EXU/ALU/_adder_io_result [29] ) );
BUF_X1 \EXU/ALU/adder/_768_ ( .A(\EXU/casez_tmp_0 [30] ), .Z(\EXU/ALU/adder/_057_ ) );
BUF_X1 \EXU/ALU/adder/_769_ ( .A(\EXU/_0023_ ), .Z(\EXU/ALU/adder/_025_ ) );
BUF_X1 \EXU/ALU/adder/_770_ ( .A(\EXU/ALU/adder/_090_ ), .Z(\EXU/ALU/_adder_io_result [30] ) );
BUF_X1 \EXU/ALU/adder/_771_ ( .A(\EXU/casez_tmp_0 [31] ), .Z(\EXU/ALU/adder/_058_ ) );
BUF_X1 \EXU/ALU/adder/_772_ ( .A(\EXU/_0024_ ), .Z(\EXU/ALU/adder/_026_ ) );
BUF_X1 \EXU/ALU/adder/_773_ ( .A(\EXU/ALU/adder/_091_ ), .Z(\EXU/ALU/_adder_io_result [31] ) );
BUF_X1 \EXU/ALU/adder/_774_ ( .A(\EXU/ALU/adder/_099_ ), .Z(\EXU/_ALU_io_zero ) );
BUF_X1 \EXU/ALU/adder/_775_ ( .A(\EXU/ALU/adder/_066_ ), .Z(\EXU/ALU/_adder_io_overflow ) );
BUF_X1 \EXU/ALU/adder/_776_ ( .A(\EXU/ALU/adder/_001_ ), .Z(\EXU/ALU/_adder_io_carry ) );
OR2_X4 \EXU/ALU/aluControl/_05_ ( .A1(\EXU/ALU/aluControl/_02_ ), .A2(\EXU/ALU/aluControl/_00_ ), .ZN(\EXU/ALU/aluControl/_04_ ) );
INV_X1 \EXU/ALU/aluControl/_06_ ( .A(\EXU/ALU/aluControl/_01_ ), .ZN(\EXU/ALU/aluControl/_03_ ) );
BUF_X1 \EXU/ALU/aluControl/_07_ ( .A(\EXU/in_control_aluCtr [0] ), .Z(\EXU/ALU/_aluControl_io_aluSel [0] ) );
BUF_X1 \EXU/ALU/aluControl/_08_ ( .A(\EXU/in_control_aluCtr [1] ), .Z(\EXU/ALU/_aluControl_io_aluSel [1] ) );
BUF_X1 \EXU/ALU/aluControl/_09_ ( .A(\EXU/in_control_aluCtr [2] ), .Z(\EXU/ALU/_aluControl_io_aluSel [2] ) );
BUF_X1 \EXU/ALU/aluControl/_10_ ( .A(\EXU/in_control_aluCtr [3] ), .Z(\EXU/ALU/_aluControl_io_isArith ) );
BUF_X1 \EXU/ALU/aluControl/_11_ ( .A(\EXU/in_control_aluCtr [3] ), .Z(\EXU/ALU/_aluControl_io_isUnsigned ) );
BUF_X1 \EXU/ALU/aluControl/_12_ ( .A(\EXU/in_control_aluCtr [3] ), .Z(\EXU/ALU/aluControl/_02_ ) );
BUF_X1 \EXU/ALU/aluControl/_13_ ( .A(\EXU/in_control_aluCtr [1] ), .Z(\EXU/ALU/aluControl/_00_ ) );
BUF_X1 \EXU/ALU/aluControl/_14_ ( .A(\EXU/ALU/aluControl/_04_ ), .Z(\EXU/ALU/_aluControl_io_isSub ) );
BUF_X1 \EXU/ALU/aluControl/_15_ ( .A(\EXU/in_control_aluCtr [2] ), .Z(\EXU/ALU/aluControl/_01_ ) );
BUF_X1 \EXU/ALU/aluControl/_16_ ( .A(\EXU/ALU/aluControl/_03_ ), .Z(\EXU/ALU/_aluControl_io_isLeft ) );
AND2_X1 \EXU/ALU/barrelShift/_0564_ ( .A1(\EXU/ALU/barrelShift/_0065_ ), .A2(\EXU/ALU/barrelShift/_0067_ ), .ZN(\EXU/ALU/barrelShift/_0536_ ) );
AND2_X4 \EXU/ALU/barrelShift/_0565_ ( .A1(\EXU/ALU/barrelShift/_0056_ ), .A2(\EXU/ALU/barrelShift/_0064_ ), .ZN(\EXU/ALU/barrelShift/_0537_ ) );
INV_X1 \EXU/ALU/barrelShift/_0566_ ( .A(\EXU/ALU/barrelShift/_0067_ ), .ZN(\EXU/ALU/barrelShift/_0538_ ) );
NOR2_X2 \EXU/ALU/barrelShift/_0567_ ( .A1(\EXU/ALU/barrelShift/_0538_ ), .A2(\EXU/ALU/barrelShift/_0065_ ), .ZN(\EXU/ALU/barrelShift/_0539_ ) );
AOI21_X1 \EXU/ALU/barrelShift/_0568_ ( .A(\EXU/ALU/barrelShift/_0065_ ), .B1(\EXU/ALU/barrelShift/_0056_ ), .B2(\EXU/ALU/barrelShift/_0064_ ), .ZN(\EXU/ALU/barrelShift/_0540_ ) );
INV_X32 \EXU/ALU/barrelShift/_0569_ ( .A(\EXU/ALU/barrelShift/_0069_ ), .ZN(\EXU/ALU/barrelShift/_0541_ ) );
NOR2_X1 \EXU/ALU/barrelShift/_0570_ ( .A1(\EXU/ALU/barrelShift/_0540_ ), .A2(\EXU/ALU/barrelShift/_0541_ ), .ZN(\EXU/ALU/barrelShift/_0542_ ) );
INV_X4 \EXU/ALU/barrelShift/_0571_ ( .A(\EXU/ALU/barrelShift/_0537_ ), .ZN(\EXU/ALU/barrelShift/_0543_ ) );
INV_X32 \EXU/ALU/barrelShift/_0572_ ( .A(\EXU/ALU/barrelShift/_0070_ ), .ZN(\EXU/ALU/barrelShift/_0544_ ) );
NOR2_X4 \EXU/ALU/barrelShift/_0573_ ( .A1(\EXU/ALU/barrelShift/_0544_ ), .A2(\EXU/ALU/barrelShift/_0065_ ), .ZN(\EXU/ALU/barrelShift/_0545_ ) );
AND2_X4 \EXU/ALU/barrelShift/_0574_ ( .A1(\EXU/ALU/barrelShift/_0543_ ), .A2(\EXU/ALU/barrelShift/_0545_ ), .ZN(\EXU/ALU/barrelShift/_0546_ ) );
BUF_X16 \EXU/ALU/barrelShift/_0575_ ( .A(\EXU/ALU/barrelShift/_0546_ ), .Z(\EXU/ALU/barrelShift/_0547_ ) );
AND2_X4 \EXU/ALU/barrelShift/_0576_ ( .A1(\EXU/ALU/barrelShift/_0070_ ), .A2(\EXU/ALU/barrelShift/_0065_ ), .ZN(\EXU/ALU/barrelShift/_0548_ ) );
INV_X4 \EXU/ALU/barrelShift/_0577_ ( .A(\EXU/ALU/barrelShift/_0548_ ), .ZN(\EXU/ALU/barrelShift/_0549_ ) );
BUF_X8 \EXU/ALU/barrelShift/_0578_ ( .A(\EXU/ALU/barrelShift/_0549_ ), .Z(\EXU/ALU/barrelShift/_0550_ ) );
NOR2_X1 \EXU/ALU/barrelShift/_0579_ ( .A1(\EXU/ALU/barrelShift/_0550_ ), .A2(\EXU/ALU/barrelShift/_0033_ ), .ZN(\EXU/ALU/barrelShift/_0551_ ) );
NOR2_X1 \EXU/ALU/barrelShift/_0580_ ( .A1(\EXU/ALU/barrelShift/_0070_ ), .A2(\EXU/ALU/barrelShift/_0050_ ), .ZN(\EXU/ALU/barrelShift/_0552_ ) );
NOR3_X4 \EXU/ALU/barrelShift/_0581_ ( .A1(\EXU/ALU/barrelShift/_0547_ ), .A2(\EXU/ALU/barrelShift/_0551_ ), .A3(\EXU/ALU/barrelShift/_0552_ ), .ZN(\EXU/ALU/barrelShift/_0553_ ) );
BUF_X2 \EXU/ALU/barrelShift/_0582_ ( .A(\EXU/ALU/barrelShift/_0541_ ), .Z(\EXU/ALU/barrelShift/_0554_ ) );
AOI21_X2 \EXU/ALU/barrelShift/_0583_ ( .A(\EXU/ALU/barrelShift/_0542_ ), .B1(\EXU/ALU/barrelShift/_0553_ ), .B2(\EXU/ALU/barrelShift/_0554_ ), .ZN(\EXU/ALU/barrelShift/_0555_ ) );
OAI22_X1 \EXU/ALU/barrelShift/_0584_ ( .A1(\EXU/ALU/barrelShift/_0549_ ), .A2(\EXU/ALU/barrelShift/_0054_ ), .B1(\EXU/ALU/barrelShift/_0070_ ), .B2(\EXU/ALU/barrelShift/_0041_ ), .ZN(\EXU/ALU/barrelShift/_0556_ ) );
NOR2_X1 \EXU/ALU/barrelShift/_0585_ ( .A1(\EXU/ALU/barrelShift/_0556_ ), .A2(\EXU/ALU/barrelShift/_0546_ ), .ZN(\EXU/ALU/barrelShift/_0557_ ) );
AND2_X2 \EXU/ALU/barrelShift/_0586_ ( .A1(\EXU/ALU/barrelShift/_0065_ ), .A2(\EXU/ALU/barrelShift/_0069_ ), .ZN(\EXU/ALU/barrelShift/_0558_ ) );
INV_X1 \EXU/ALU/barrelShift/_0587_ ( .A(\EXU/ALU/barrelShift/_0558_ ), .ZN(\EXU/ALU/barrelShift/_0559_ ) );
BUF_X4 \EXU/ALU/barrelShift/_0588_ ( .A(\EXU/ALU/barrelShift/_0559_ ), .Z(\EXU/ALU/barrelShift/_0560_ ) );
NOR2_X1 \EXU/ALU/barrelShift/_0589_ ( .A1(\EXU/ALU/barrelShift/_0557_ ), .A2(\EXU/ALU/barrelShift/_0560_ ), .ZN(\EXU/ALU/barrelShift/_0561_ ) );
NOR2_X4 \EXU/ALU/barrelShift/_0590_ ( .A1(\EXU/ALU/barrelShift/_0555_ ), .A2(\EXU/ALU/barrelShift/_0561_ ), .ZN(\EXU/ALU/barrelShift/_0562_ ) );
OAI22_X2 \EXU/ALU/barrelShift/_0591_ ( .A1(\EXU/ALU/barrelShift/_0550_ ), .A2(\EXU/ALU/barrelShift/_0060_ ), .B1(\EXU/ALU/barrelShift/_0070_ ), .B2(\EXU/ALU/barrelShift/_0046_ ), .ZN(\EXU/ALU/barrelShift/_0563_ ) );
OAI21_X2 \EXU/ALU/barrelShift/_0592_ ( .A(\EXU/ALU/barrelShift/_0558_ ), .B1(\EXU/ALU/barrelShift/_0563_ ), .B2(\EXU/ALU/barrelShift/_0547_ ), .ZN(\EXU/ALU/barrelShift/_0071_ ) );
NOR2_X1 \EXU/ALU/barrelShift/_0593_ ( .A1(\EXU/ALU/barrelShift/_0549_ ), .A2(\EXU/ALU/barrelShift/_0037_ ), .ZN(\EXU/ALU/barrelShift/_0072_ ) );
NOR2_X1 \EXU/ALU/barrelShift/_0594_ ( .A1(\EXU/ALU/barrelShift/_0070_ ), .A2(\EXU/ALU/barrelShift/_0055_ ), .ZN(\EXU/ALU/barrelShift/_0073_ ) );
NOR3_X2 \EXU/ALU/barrelShift/_0595_ ( .A1(\EXU/ALU/barrelShift/_0546_ ), .A2(\EXU/ALU/barrelShift/_0072_ ), .A3(\EXU/ALU/barrelShift/_0073_ ), .ZN(\EXU/ALU/barrelShift/_0074_ ) );
AND2_X1 \EXU/ALU/barrelShift/_0596_ ( .A1(\EXU/ALU/barrelShift/_0074_ ), .A2(\EXU/ALU/barrelShift/_0554_ ), .ZN(\EXU/ALU/barrelShift/_0075_ ) );
OAI21_X1 \EXU/ALU/barrelShift/_0597_ ( .A(\EXU/ALU/barrelShift/_0071_ ), .B1(\EXU/ALU/barrelShift/_0075_ ), .B2(\EXU/ALU/barrelShift/_0542_ ), .ZN(\EXU/ALU/barrelShift/_0076_ ) );
INV_X2 \EXU/ALU/barrelShift/_0598_ ( .A(\EXU/ALU/barrelShift/_0068_ ), .ZN(\EXU/ALU/barrelShift/_0077_ ) );
NOR2_X1 \EXU/ALU/barrelShift/_0599_ ( .A1(\EXU/ALU/barrelShift/_0077_ ), .A2(\EXU/ALU/barrelShift/_0065_ ), .ZN(\EXU/ALU/barrelShift/_0078_ ) );
INV_X2 \EXU/ALU/barrelShift/_0600_ ( .A(\EXU/ALU/barrelShift/_0078_ ), .ZN(\EXU/ALU/barrelShift/_0079_ ) );
OAI22_X1 \EXU/ALU/barrelShift/_0601_ ( .A1(\EXU/ALU/barrelShift/_0076_ ), .A2(\EXU/ALU/barrelShift/_0068_ ), .B1(\EXU/ALU/barrelShift/_0543_ ), .B2(\EXU/ALU/barrelShift/_0079_ ), .ZN(\EXU/ALU/barrelShift/_0080_ ) );
AND2_X2 \EXU/ALU/barrelShift/_0602_ ( .A1(\EXU/ALU/barrelShift/_0065_ ), .A2(\EXU/ALU/barrelShift/_0068_ ), .ZN(\EXU/ALU/barrelShift/_0081_ ) );
INV_X1 \EXU/ALU/barrelShift/_0603_ ( .A(\EXU/ALU/barrelShift/_0081_ ), .ZN(\EXU/ALU/barrelShift/_0082_ ) );
BUF_X4 \EXU/ALU/barrelShift/_0604_ ( .A(\EXU/ALU/barrelShift/_0082_ ), .Z(\EXU/ALU/barrelShift/_0083_ ) );
MUX2_X2 \EXU/ALU/barrelShift/_0605_ ( .A(\EXU/ALU/barrelShift/_0562_ ), .B(\EXU/ALU/barrelShift/_0080_ ), .S(\EXU/ALU/barrelShift/_0083_ ), .Z(\EXU/ALU/barrelShift/_0084_ ) );
AOI221_X2 \EXU/ALU/barrelShift/_0606_ ( .A(\EXU/ALU/barrelShift/_0536_ ), .B1(\EXU/ALU/barrelShift/_0537_ ), .B2(\EXU/ALU/barrelShift/_0539_ ), .C1(\EXU/ALU/barrelShift/_0084_ ), .C2(\EXU/ALU/barrelShift/_0538_ ), .ZN(\EXU/ALU/barrelShift/_0085_ ) );
BUF_X4 \EXU/ALU/barrelShift/_0607_ ( .A(\EXU/ALU/barrelShift/_0536_ ), .Z(\EXU/ALU/barrelShift/_0086_ ) );
BUF_X4 \EXU/ALU/barrelShift/_0608_ ( .A(\EXU/ALU/barrelShift/_0086_ ), .Z(\EXU/ALU/barrelShift/_0087_ ) );
OAI22_X1 \EXU/ALU/barrelShift/_0609_ ( .A1(\EXU/ALU/barrelShift/_0550_ ), .A2(\EXU/ALU/barrelShift/_0058_ ), .B1(\EXU/ALU/barrelShift/_0070_ ), .B2(\EXU/ALU/barrelShift/_0044_ ), .ZN(\EXU/ALU/barrelShift/_0088_ ) );
NOR2_X4 \EXU/ALU/barrelShift/_0610_ ( .A1(\EXU/ALU/barrelShift/_0088_ ), .A2(\EXU/ALU/barrelShift/_0547_ ), .ZN(\EXU/ALU/barrelShift/_0089_ ) );
NOR2_X2 \EXU/ALU/barrelShift/_0611_ ( .A1(\EXU/ALU/barrelShift/_0089_ ), .A2(\EXU/ALU/barrelShift/_0560_ ), .ZN(\EXU/ALU/barrelShift/_0090_ ) );
INV_X1 \EXU/ALU/barrelShift/_0612_ ( .A(\EXU/ALU/barrelShift/_0542_ ), .ZN(\EXU/ALU/barrelShift/_0091_ ) );
OAI22_X1 \EXU/ALU/barrelShift/_0613_ ( .A1(\EXU/ALU/barrelShift/_0550_ ), .A2(\EXU/ALU/barrelShift/_0035_ ), .B1(\EXU/ALU/barrelShift/_0070_ ), .B2(\EXU/ALU/barrelShift/_0052_ ), .ZN(\EXU/ALU/barrelShift/_0092_ ) );
NOR2_X4 \EXU/ALU/barrelShift/_0614_ ( .A1(\EXU/ALU/barrelShift/_0092_ ), .A2(\EXU/ALU/barrelShift/_0547_ ), .ZN(\EXU/ALU/barrelShift/_0093_ ) );
BUF_X4 \EXU/ALU/barrelShift/_0615_ ( .A(\EXU/ALU/barrelShift/_0541_ ), .Z(\EXU/ALU/barrelShift/_0094_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0616_ ( .A1(\EXU/ALU/barrelShift/_0093_ ), .A2(\EXU/ALU/barrelShift/_0094_ ), .ZN(\EXU/ALU/barrelShift/_0095_ ) );
AOI21_X2 \EXU/ALU/barrelShift/_0617_ ( .A(\EXU/ALU/barrelShift/_0090_ ), .B1(\EXU/ALU/barrelShift/_0091_ ), .B2(\EXU/ALU/barrelShift/_0095_ ), .ZN(\EXU/ALU/barrelShift/_0096_ ) );
BUF_X4 \EXU/ALU/barrelShift/_0618_ ( .A(\EXU/ALU/barrelShift/_0077_ ), .Z(\EXU/ALU/barrelShift/_0097_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0619_ ( .A1(\EXU/ALU/barrelShift/_0096_ ), .A2(\EXU/ALU/barrelShift/_0097_ ), .ZN(\EXU/ALU/barrelShift/_0098_ ) );
OR2_X1 \EXU/ALU/barrelShift/_0620_ ( .A1(\EXU/ALU/barrelShift/_0540_ ), .A2(\EXU/ALU/barrelShift/_0077_ ), .ZN(\EXU/ALU/barrelShift/_0099_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0621_ ( .A1(\EXU/ALU/barrelShift/_0098_ ), .A2(\EXU/ALU/barrelShift/_0099_ ), .ZN(\EXU/ALU/barrelShift/_0100_ ) );
BUF_X4 \EXU/ALU/barrelShift/_0622_ ( .A(\EXU/ALU/barrelShift/_0081_ ), .Z(\EXU/ALU/barrelShift/_0101_ ) );
OAI22_X2 \EXU/ALU/barrelShift/_0623_ ( .A1(\EXU/ALU/barrelShift/_0550_ ), .A2(\EXU/ALU/barrelShift/_0062_ ), .B1(\EXU/ALU/barrelShift/_0070_ ), .B2(\EXU/ALU/barrelShift/_0048_ ), .ZN(\EXU/ALU/barrelShift/_0102_ ) );
NOR2_X2 \EXU/ALU/barrelShift/_0624_ ( .A1(\EXU/ALU/barrelShift/_0102_ ), .A2(\EXU/ALU/barrelShift/_0546_ ), .ZN(\EXU/ALU/barrelShift/_0103_ ) );
AOI21_X1 \EXU/ALU/barrelShift/_0625_ ( .A(\EXU/ALU/barrelShift/_0542_ ), .B1(\EXU/ALU/barrelShift/_0103_ ), .B2(\EXU/ALU/barrelShift/_0554_ ), .ZN(\EXU/ALU/barrelShift/_0104_ ) );
OAI22_X1 \EXU/ALU/barrelShift/_0626_ ( .A1(\EXU/ALU/barrelShift/_0549_ ), .A2(\EXU/ALU/barrelShift/_0032_ ), .B1(\EXU/ALU/barrelShift/_0070_ ), .B2(\EXU/ALU/barrelShift/_0039_ ), .ZN(\EXU/ALU/barrelShift/_0105_ ) );
NOR2_X2 \EXU/ALU/barrelShift/_0627_ ( .A1(\EXU/ALU/barrelShift/_0105_ ), .A2(\EXU/ALU/barrelShift/_0546_ ), .ZN(\EXU/ALU/barrelShift/_0106_ ) );
NOR2_X1 \EXU/ALU/barrelShift/_0628_ ( .A1(\EXU/ALU/barrelShift/_0106_ ), .A2(\EXU/ALU/barrelShift/_0559_ ), .ZN(\EXU/ALU/barrelShift/_0107_ ) );
OAI21_X1 \EXU/ALU/barrelShift/_0629_ ( .A(\EXU/ALU/barrelShift/_0101_ ), .B1(\EXU/ALU/barrelShift/_0104_ ), .B2(\EXU/ALU/barrelShift/_0107_ ), .ZN(\EXU/ALU/barrelShift/_0108_ ) );
NAND2_X2 \EXU/ALU/barrelShift/_0630_ ( .A1(\EXU/ALU/barrelShift/_0100_ ), .A2(\EXU/ALU/barrelShift/_0108_ ), .ZN(\EXU/ALU/barrelShift/_0109_ ) );
AOI21_X2 \EXU/ALU/barrelShift/_0631_ ( .A(\EXU/ALU/barrelShift/_0085_ ), .B1(\EXU/ALU/barrelShift/_0087_ ), .B2(\EXU/ALU/barrelShift/_0109_ ), .ZN(\EXU/ALU/barrelShift/_0110_ ) );
INV_X1 \EXU/ALU/barrelShift/_0632_ ( .A(\EXU/ALU/barrelShift/_0066_ ), .ZN(\EXU/ALU/barrelShift/_0111_ ) );
BUF_X4 \EXU/ALU/barrelShift/_0633_ ( .A(\EXU/ALU/barrelShift/_0111_ ), .Z(\EXU/ALU/barrelShift/_0112_ ) );
BUF_X4 \EXU/ALU/barrelShift/_0634_ ( .A(\EXU/ALU/barrelShift/_0112_ ), .Z(\EXU/ALU/barrelShift/_0113_ ) );
AND2_X1 \EXU/ALU/barrelShift/_0635_ ( .A1(\EXU/ALU/barrelShift/_0065_ ), .A2(\EXU/ALU/barrelShift/_0066_ ), .ZN(\EXU/ALU/barrelShift/_0114_ ) );
BUF_X4 \EXU/ALU/barrelShift/_0636_ ( .A(\EXU/ALU/barrelShift/_0114_ ), .Z(\EXU/ALU/barrelShift/_0115_ ) );
OAI22_X2 \EXU/ALU/barrelShift/_0637_ ( .A1(\EXU/ALU/barrelShift/_0550_ ), .A2(\EXU/ALU/barrelShift/_0034_ ), .B1(\EXU/ALU/barrelShift/_0070_ ), .B2(\EXU/ALU/barrelShift/_0051_ ), .ZN(\EXU/ALU/barrelShift/_0116_ ) );
NOR2_X4 \EXU/ALU/barrelShift/_0638_ ( .A1(\EXU/ALU/barrelShift/_0116_ ), .A2(\EXU/ALU/barrelShift/_0547_ ), .ZN(\EXU/ALU/barrelShift/_0117_ ) );
AOI21_X2 \EXU/ALU/barrelShift/_0639_ ( .A(\EXU/ALU/barrelShift/_0542_ ), .B1(\EXU/ALU/barrelShift/_0117_ ), .B2(\EXU/ALU/barrelShift/_0554_ ), .ZN(\EXU/ALU/barrelShift/_0118_ ) );
OAI22_X1 \EXU/ALU/barrelShift/_0640_ ( .A1(\EXU/ALU/barrelShift/_0550_ ), .A2(\EXU/ALU/barrelShift/_0057_ ), .B1(\EXU/ALU/barrelShift/_0070_ ), .B2(\EXU/ALU/barrelShift/_0042_ ), .ZN(\EXU/ALU/barrelShift/_0119_ ) );
NOR2_X4 \EXU/ALU/barrelShift/_0641_ ( .A1(\EXU/ALU/barrelShift/_0119_ ), .A2(\EXU/ALU/barrelShift/_0547_ ), .ZN(\EXU/ALU/barrelShift/_0120_ ) );
NOR2_X2 \EXU/ALU/barrelShift/_0642_ ( .A1(\EXU/ALU/barrelShift/_0120_ ), .A2(\EXU/ALU/barrelShift/_0560_ ), .ZN(\EXU/ALU/barrelShift/_0121_ ) );
NOR2_X2 \EXU/ALU/barrelShift/_0643_ ( .A1(\EXU/ALU/barrelShift/_0118_ ), .A2(\EXU/ALU/barrelShift/_0121_ ), .ZN(\EXU/ALU/barrelShift/_0122_ ) );
BUF_X2 \EXU/ALU/barrelShift/_0644_ ( .A(\EXU/ALU/barrelShift/_0558_ ), .Z(\EXU/ALU/barrelShift/_0123_ ) );
OAI22_X1 \EXU/ALU/barrelShift/_0645_ ( .A1(\EXU/ALU/barrelShift/_0549_ ), .A2(\EXU/ALU/barrelShift/_0061_ ), .B1(\EXU/ALU/barrelShift/_0070_ ), .B2(\EXU/ALU/barrelShift/_0047_ ), .ZN(\EXU/ALU/barrelShift/_0124_ ) );
OAI21_X2 \EXU/ALU/barrelShift/_0646_ ( .A(\EXU/ALU/barrelShift/_0123_ ), .B1(\EXU/ALU/barrelShift/_0124_ ), .B2(\EXU/ALU/barrelShift/_0547_ ), .ZN(\EXU/ALU/barrelShift/_0125_ ) );
AND2_X2 \EXU/ALU/barrelShift/_0647_ ( .A1(\EXU/ALU/barrelShift/_0545_ ), .A2(\EXU/ALU/barrelShift/_0537_ ), .ZN(\EXU/ALU/barrelShift/_0126_ ) );
AOI21_X1 \EXU/ALU/barrelShift/_0648_ ( .A(\EXU/ALU/barrelShift/_0126_ ), .B1(\EXU/ALU/barrelShift/_0544_ ), .B2(\EXU/ALU/barrelShift/_0056_ ), .ZN(\EXU/ALU/barrelShift/_0127_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0649_ ( .A1(\EXU/ALU/barrelShift/_0070_ ), .A2(\EXU/ALU/barrelShift/_0065_ ), .A3(\EXU/ALU/barrelShift/_0038_ ), .ZN(\EXU/ALU/barrelShift/_0128_ ) );
AOI21_X1 \EXU/ALU/barrelShift/_0650_ ( .A(\EXU/ALU/barrelShift/_0069_ ), .B1(\EXU/ALU/barrelShift/_0127_ ), .B2(\EXU/ALU/barrelShift/_0128_ ), .ZN(\EXU/ALU/barrelShift/_0129_ ) );
OAI21_X1 \EXU/ALU/barrelShift/_0651_ ( .A(\EXU/ALU/barrelShift/_0125_ ), .B1(\EXU/ALU/barrelShift/_0129_ ), .B2(\EXU/ALU/barrelShift/_0542_ ), .ZN(\EXU/ALU/barrelShift/_0130_ ) );
OAI22_X1 \EXU/ALU/barrelShift/_0652_ ( .A1(\EXU/ALU/barrelShift/_0130_ ), .A2(\EXU/ALU/barrelShift/_0068_ ), .B1(\EXU/ALU/barrelShift/_0543_ ), .B2(\EXU/ALU/barrelShift/_0079_ ), .ZN(\EXU/ALU/barrelShift/_0131_ ) );
BUF_X4 \EXU/ALU/barrelShift/_0653_ ( .A(\EXU/ALU/barrelShift/_0083_ ), .Z(\EXU/ALU/barrelShift/_0132_ ) );
MUX2_X2 \EXU/ALU/barrelShift/_0654_ ( .A(\EXU/ALU/barrelShift/_0122_ ), .B(\EXU/ALU/barrelShift/_0131_ ), .S(\EXU/ALU/barrelShift/_0132_ ), .Z(\EXU/ALU/barrelShift/_0133_ ) );
OAI22_X1 \EXU/ALU/barrelShift/_0655_ ( .A1(\EXU/ALU/barrelShift/_0550_ ), .A2(\EXU/ALU/barrelShift/_0059_ ), .B1(\EXU/ALU/barrelShift/_0070_ ), .B2(\EXU/ALU/barrelShift/_0045_ ), .ZN(\EXU/ALU/barrelShift/_0134_ ) );
NOR2_X4 \EXU/ALU/barrelShift/_0656_ ( .A1(\EXU/ALU/barrelShift/_0134_ ), .A2(\EXU/ALU/barrelShift/_0547_ ), .ZN(\EXU/ALU/barrelShift/_0135_ ) );
NOR2_X2 \EXU/ALU/barrelShift/_0657_ ( .A1(\EXU/ALU/barrelShift/_0135_ ), .A2(\EXU/ALU/barrelShift/_0560_ ), .ZN(\EXU/ALU/barrelShift/_0136_ ) );
OAI22_X1 \EXU/ALU/barrelShift/_0658_ ( .A1(\EXU/ALU/barrelShift/_0550_ ), .A2(\EXU/ALU/barrelShift/_0036_ ), .B1(\EXU/ALU/barrelShift/_0070_ ), .B2(\EXU/ALU/barrelShift/_0053_ ), .ZN(\EXU/ALU/barrelShift/_0137_ ) );
NOR2_X4 \EXU/ALU/barrelShift/_0659_ ( .A1(\EXU/ALU/barrelShift/_0137_ ), .A2(\EXU/ALU/barrelShift/_0547_ ), .ZN(\EXU/ALU/barrelShift/_0138_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0660_ ( .A1(\EXU/ALU/barrelShift/_0138_ ), .A2(\EXU/ALU/barrelShift/_0554_ ), .ZN(\EXU/ALU/barrelShift/_0139_ ) );
AOI21_X2 \EXU/ALU/barrelShift/_0661_ ( .A(\EXU/ALU/barrelShift/_0136_ ), .B1(\EXU/ALU/barrelShift/_0091_ ), .B2(\EXU/ALU/barrelShift/_0139_ ), .ZN(\EXU/ALU/barrelShift/_0140_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0662_ ( .A1(\EXU/ALU/barrelShift/_0140_ ), .A2(\EXU/ALU/barrelShift/_0097_ ), .ZN(\EXU/ALU/barrelShift/_0141_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0663_ ( .A1(\EXU/ALU/barrelShift/_0141_ ), .A2(\EXU/ALU/barrelShift/_0099_ ), .ZN(\EXU/ALU/barrelShift/_0142_ ) );
OAI22_X1 \EXU/ALU/barrelShift/_0664_ ( .A1(\EXU/ALU/barrelShift/_0550_ ), .A2(\EXU/ALU/barrelShift/_0063_ ), .B1(\EXU/ALU/barrelShift/_0070_ ), .B2(\EXU/ALU/barrelShift/_0049_ ), .ZN(\EXU/ALU/barrelShift/_0143_ ) );
NOR2_X1 \EXU/ALU/barrelShift/_0665_ ( .A1(\EXU/ALU/barrelShift/_0143_ ), .A2(\EXU/ALU/barrelShift/_0546_ ), .ZN(\EXU/ALU/barrelShift/_0144_ ) );
AOI21_X1 \EXU/ALU/barrelShift/_0666_ ( .A(\EXU/ALU/barrelShift/_0542_ ), .B1(\EXU/ALU/barrelShift/_0144_ ), .B2(\EXU/ALU/barrelShift/_0554_ ), .ZN(\EXU/ALU/barrelShift/_0145_ ) );
OAI22_X1 \EXU/ALU/barrelShift/_0667_ ( .A1(\EXU/ALU/barrelShift/_0549_ ), .A2(\EXU/ALU/barrelShift/_0043_ ), .B1(\EXU/ALU/barrelShift/_0070_ ), .B2(\EXU/ALU/barrelShift/_0040_ ), .ZN(\EXU/ALU/barrelShift/_0146_ ) );
NOR2_X2 \EXU/ALU/barrelShift/_0668_ ( .A1(\EXU/ALU/barrelShift/_0146_ ), .A2(\EXU/ALU/barrelShift/_0546_ ), .ZN(\EXU/ALU/barrelShift/_0147_ ) );
NOR2_X1 \EXU/ALU/barrelShift/_0669_ ( .A1(\EXU/ALU/barrelShift/_0147_ ), .A2(\EXU/ALU/barrelShift/_0559_ ), .ZN(\EXU/ALU/barrelShift/_0148_ ) );
OAI21_X1 \EXU/ALU/barrelShift/_0670_ ( .A(\EXU/ALU/barrelShift/_0101_ ), .B1(\EXU/ALU/barrelShift/_0145_ ), .B2(\EXU/ALU/barrelShift/_0148_ ), .ZN(\EXU/ALU/barrelShift/_0149_ ) );
AND2_X2 \EXU/ALU/barrelShift/_0671_ ( .A1(\EXU/ALU/barrelShift/_0142_ ), .A2(\EXU/ALU/barrelShift/_0149_ ), .ZN(\EXU/ALU/barrelShift/_0150_ ) );
BUF_X4 \EXU/ALU/barrelShift/_0672_ ( .A(\EXU/ALU/barrelShift/_0538_ ), .Z(\EXU/ALU/barrelShift/_0151_ ) );
AOI22_X2 \EXU/ALU/barrelShift/_0673_ ( .A1(\EXU/ALU/barrelShift/_0133_ ), .A2(\EXU/ALU/barrelShift/_0539_ ), .B1(\EXU/ALU/barrelShift/_0150_ ), .B2(\EXU/ALU/barrelShift/_0151_ ), .ZN(\EXU/ALU/barrelShift/_0152_ ) );
INV_X1 \EXU/ALU/barrelShift/_0674_ ( .A(\EXU/ALU/barrelShift/_0086_ ), .ZN(\EXU/ALU/barrelShift/_0153_ ) );
NOR2_X2 \EXU/ALU/barrelShift/_0675_ ( .A1(\EXU/ALU/barrelShift/_0124_ ), .A2(\EXU/ALU/barrelShift/_0546_ ), .ZN(\EXU/ALU/barrelShift/_0154_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0676_ ( .A1(\EXU/ALU/barrelShift/_0545_ ), .A2(\EXU/ALU/barrelShift/_0056_ ), .ZN(\EXU/ALU/barrelShift/_0155_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0677_ ( .A1(\EXU/ALU/barrelShift/_0544_ ), .A2(\EXU/ALU/barrelShift/_0038_ ), .ZN(\EXU/ALU/barrelShift/_0156_ ) );
AND2_X1 \EXU/ALU/barrelShift/_0678_ ( .A1(\EXU/ALU/barrelShift/_0155_ ), .A2(\EXU/ALU/barrelShift/_0156_ ), .ZN(\EXU/ALU/barrelShift/_0157_ ) );
INV_X1 \EXU/ALU/barrelShift/_0679_ ( .A(\EXU/ALU/barrelShift/_0157_ ), .ZN(\EXU/ALU/barrelShift/_0158_ ) );
AOI22_X1 \EXU/ALU/barrelShift/_0680_ ( .A1(\EXU/ALU/barrelShift/_0554_ ), .A2(\EXU/ALU/barrelShift/_0154_ ), .B1(\EXU/ALU/barrelShift/_0158_ ), .B2(\EXU/ALU/barrelShift/_0558_ ), .ZN(\EXU/ALU/barrelShift/_0159_ ) );
INV_X1 \EXU/ALU/barrelShift/_0681_ ( .A(\EXU/ALU/barrelShift/_0159_ ), .ZN(\EXU/ALU/barrelShift/_0160_ ) );
NOR2_X4 \EXU/ALU/barrelShift/_0682_ ( .A1(\EXU/ALU/barrelShift/_0541_ ), .A2(\EXU/ALU/barrelShift/_0065_ ), .ZN(\EXU/ALU/barrelShift/_0161_ ) );
INV_X1 \EXU/ALU/barrelShift/_0683_ ( .A(\EXU/ALU/barrelShift/_0161_ ), .ZN(\EXU/ALU/barrelShift/_0162_ ) );
BUF_X4 \EXU/ALU/barrelShift/_0684_ ( .A(\EXU/ALU/barrelShift/_0162_ ), .Z(\EXU/ALU/barrelShift/_0163_ ) );
AOI21_X1 \EXU/ALU/barrelShift/_0685_ ( .A(\EXU/ALU/barrelShift/_0163_ ), .B1(\EXU/ALU/barrelShift/_0127_ ), .B2(\EXU/ALU/barrelShift/_0128_ ), .ZN(\EXU/ALU/barrelShift/_0164_ ) );
NOR2_X1 \EXU/ALU/barrelShift/_0686_ ( .A1(\EXU/ALU/barrelShift/_0160_ ), .A2(\EXU/ALU/barrelShift/_0164_ ), .ZN(\EXU/ALU/barrelShift/_0165_ ) );
INV_X1 \EXU/ALU/barrelShift/_0687_ ( .A(\EXU/ALU/barrelShift/_0165_ ), .ZN(\EXU/ALU/barrelShift/_0166_ ) );
AOI22_X1 \EXU/ALU/barrelShift/_0688_ ( .A1(\EXU/ALU/barrelShift/_0166_ ), .A2(\EXU/ALU/barrelShift/_0101_ ), .B1(\EXU/ALU/barrelShift/_0097_ ), .B2(\EXU/ALU/barrelShift/_0122_ ), .ZN(\EXU/ALU/barrelShift/_0167_ ) );
OR2_X1 \EXU/ALU/barrelShift/_0689_ ( .A1(\EXU/ALU/barrelShift/_0130_ ), .A2(\EXU/ALU/barrelShift/_0079_ ), .ZN(\EXU/ALU/barrelShift/_0168_ ) );
AND2_X1 \EXU/ALU/barrelShift/_0690_ ( .A1(\EXU/ALU/barrelShift/_0167_ ), .A2(\EXU/ALU/barrelShift/_0168_ ), .ZN(\EXU/ALU/barrelShift/_0169_ ) );
OAI21_X1 \EXU/ALU/barrelShift/_0691_ ( .A(\EXU/ALU/barrelShift/_0152_ ), .B1(\EXU/ALU/barrelShift/_0153_ ), .B2(\EXU/ALU/barrelShift/_0169_ ), .ZN(\EXU/ALU/barrelShift/_0170_ ) );
AOI22_X1 \EXU/ALU/barrelShift/_0692_ ( .A1(\EXU/ALU/barrelShift/_0110_ ), .A2(\EXU/ALU/barrelShift/_0113_ ), .B1(\EXU/ALU/barrelShift/_0115_ ), .B2(\EXU/ALU/barrelShift/_0170_ ), .ZN(\EXU/ALU/barrelShift/_0171_ ) );
AOI21_X1 \EXU/ALU/barrelShift/_0693_ ( .A(\EXU/ALU/barrelShift/_0153_ ), .B1(\EXU/ALU/barrelShift/_0142_ ), .B2(\EXU/ALU/barrelShift/_0149_ ), .ZN(\EXU/ALU/barrelShift/_0172_ ) );
AOI22_X1 \EXU/ALU/barrelShift/_0694_ ( .A1(\EXU/ALU/barrelShift/_0133_ ), .A2(\EXU/ALU/barrelShift/_0151_ ), .B1(\EXU/ALU/barrelShift/_0537_ ), .B2(\EXU/ALU/barrelShift/_0539_ ), .ZN(\EXU/ALU/barrelShift/_0173_ ) );
BUF_X4 \EXU/ALU/barrelShift/_0695_ ( .A(\EXU/ALU/barrelShift/_0153_ ), .Z(\EXU/ALU/barrelShift/_0174_ ) );
AOI21_X1 \EXU/ALU/barrelShift/_0696_ ( .A(\EXU/ALU/barrelShift/_0172_ ), .B1(\EXU/ALU/barrelShift/_0173_ ), .B2(\EXU/ALU/barrelShift/_0174_ ), .ZN(\EXU/ALU/barrelShift/_0175_ ) );
NOR2_X1 \EXU/ALU/barrelShift/_0697_ ( .A1(\EXU/ALU/barrelShift/_0111_ ), .A2(\EXU/ALU/barrelShift/_0065_ ), .ZN(\EXU/ALU/barrelShift/_0176_ ) );
BUF_X4 \EXU/ALU/barrelShift/_0698_ ( .A(\EXU/ALU/barrelShift/_0176_ ), .Z(\EXU/ALU/barrelShift/_0177_ ) );
BUF_X4 \EXU/ALU/barrelShift/_0699_ ( .A(\EXU/ALU/barrelShift/_0177_ ), .Z(\EXU/ALU/barrelShift/_0178_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0700_ ( .A1(\EXU/ALU/barrelShift/_0175_ ), .A2(\EXU/ALU/barrelShift/_0178_ ), .ZN(\EXU/ALU/barrelShift/_0179_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0701_ ( .A1(\EXU/ALU/barrelShift/_0171_ ), .A2(\EXU/ALU/barrelShift/_0179_ ), .ZN(\EXU/ALU/barrelShift/_0031_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0702_ ( .A1(\EXU/ALU/barrelShift/_0110_ ), .A2(\EXU/ALU/barrelShift/_0115_ ), .ZN(\EXU/ALU/barrelShift/_0180_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0703_ ( .A1(\EXU/ALU/barrelShift/_0175_ ), .A2(\EXU/ALU/barrelShift/_0112_ ), .ZN(\EXU/ALU/barrelShift/_0181_ ) );
INV_X1 \EXU/ALU/barrelShift/_0704_ ( .A(\EXU/ALU/barrelShift/_0177_ ), .ZN(\EXU/ALU/barrelShift/_0182_ ) );
OAI211_X2 \EXU/ALU/barrelShift/_0705_ ( .A(\EXU/ALU/barrelShift/_0180_ ), .B(\EXU/ALU/barrelShift/_0181_ ), .C1(\EXU/ALU/barrelShift/_0182_ ), .C2(\EXU/ALU/barrelShift/_0543_ ), .ZN(\EXU/ALU/barrelShift/_0030_ ) );
BUF_X4 \EXU/ALU/barrelShift/_0706_ ( .A(\EXU/ALU/barrelShift/_0151_ ), .Z(\EXU/ALU/barrelShift/_0183_ ) );
NOR2_X1 \EXU/ALU/barrelShift/_0707_ ( .A1(\EXU/ALU/barrelShift/_0145_ ), .A2(\EXU/ALU/barrelShift/_0148_ ), .ZN(\EXU/ALU/barrelShift/_0184_ ) );
BUF_X2 \EXU/ALU/barrelShift/_0708_ ( .A(\EXU/ALU/barrelShift/_0078_ ), .Z(\EXU/ALU/barrelShift/_0185_ ) );
AOI221_X1 \EXU/ALU/barrelShift/_0709_ ( .A(\EXU/ALU/barrelShift/_0081_ ), .B1(\EXU/ALU/barrelShift/_0184_ ), .B2(\EXU/ALU/barrelShift/_0077_ ), .C1(\EXU/ALU/barrelShift/_0185_ ), .C2(\EXU/ALU/barrelShift/_0140_ ), .ZN(\EXU/ALU/barrelShift/_0186_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0710_ ( .A1(\EXU/ALU/barrelShift/_0545_ ), .A2(\EXU/ALU/barrelShift/_0053_ ), .ZN(\EXU/ALU/barrelShift/_0187_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0711_ ( .A1(\EXU/ALU/barrelShift/_0544_ ), .A2(\EXU/ALU/barrelShift/_0036_ ), .ZN(\EXU/ALU/barrelShift/_0188_ ) );
AND2_X1 \EXU/ALU/barrelShift/_0712_ ( .A1(\EXU/ALU/barrelShift/_0187_ ), .A2(\EXU/ALU/barrelShift/_0188_ ), .ZN(\EXU/ALU/barrelShift/_0189_ ) );
INV_X1 \EXU/ALU/barrelShift/_0713_ ( .A(\EXU/ALU/barrelShift/_0189_ ), .ZN(\EXU/ALU/barrelShift/_0190_ ) );
OAI22_X2 \EXU/ALU/barrelShift/_0714_ ( .A1(\EXU/ALU/barrelShift/_0135_ ), .A2(\EXU/ALU/barrelShift/_0069_ ), .B1(\EXU/ALU/barrelShift/_0190_ ), .B2(\EXU/ALU/barrelShift/_0560_ ), .ZN(\EXU/ALU/barrelShift/_0191_ ) );
NOR2_X1 \EXU/ALU/barrelShift/_0715_ ( .A1(\EXU/ALU/barrelShift/_0138_ ), .A2(\EXU/ALU/barrelShift/_0163_ ), .ZN(\EXU/ALU/barrelShift/_0192_ ) );
NOR2_X2 \EXU/ALU/barrelShift/_0716_ ( .A1(\EXU/ALU/barrelShift/_0191_ ), .A2(\EXU/ALU/barrelShift/_0192_ ), .ZN(\EXU/ALU/barrelShift/_0193_ ) );
NOR2_X1 \EXU/ALU/barrelShift/_0717_ ( .A1(\EXU/ALU/barrelShift/_0193_ ), .A2(\EXU/ALU/barrelShift/_0132_ ), .ZN(\EXU/ALU/barrelShift/_0194_ ) );
OR2_X2 \EXU/ALU/barrelShift/_0718_ ( .A1(\EXU/ALU/barrelShift/_0186_ ), .A2(\EXU/ALU/barrelShift/_0194_ ), .ZN(\EXU/ALU/barrelShift/_0195_ ) );
AOI22_X1 \EXU/ALU/barrelShift/_0719_ ( .A1(\EXU/ALU/barrelShift/_0183_ ), .A2(\EXU/ALU/barrelShift/_0169_ ), .B1(\EXU/ALU/barrelShift/_0195_ ), .B2(\EXU/ALU/barrelShift/_0087_ ), .ZN(\EXU/ALU/barrelShift/_0196_ ) );
BUF_X4 \EXU/ALU/barrelShift/_0720_ ( .A(\EXU/ALU/barrelShift/_0115_ ), .Z(\EXU/ALU/barrelShift/_0197_ ) );
INV_X1 \EXU/ALU/barrelShift/_0721_ ( .A(\EXU/ALU/barrelShift/_0539_ ), .ZN(\EXU/ALU/barrelShift/_0198_ ) );
BUF_X4 \EXU/ALU/barrelShift/_0722_ ( .A(\EXU/ALU/barrelShift/_0198_ ), .Z(\EXU/ALU/barrelShift/_0199_ ) );
OR2_X1 \EXU/ALU/barrelShift/_0723_ ( .A1(\EXU/ALU/barrelShift/_0150_ ), .A2(\EXU/ALU/barrelShift/_0199_ ), .ZN(\EXU/ALU/barrelShift/_0200_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0724_ ( .A1(\EXU/ALU/barrelShift/_0196_ ), .A2(\EXU/ALU/barrelShift/_0197_ ), .A3(\EXU/ALU/barrelShift/_0200_ ), .ZN(\EXU/ALU/barrelShift/_0201_ ) );
OR2_X1 \EXU/ALU/barrelShift/_0725_ ( .A1(\EXU/ALU/barrelShift/_0084_ ), .A2(\EXU/ALU/barrelShift/_0199_ ), .ZN(\EXU/ALU/barrelShift/_0202_ ) );
AND2_X1 \EXU/ALU/barrelShift/_0726_ ( .A1(\EXU/ALU/barrelShift/_0076_ ), .A2(\EXU/ALU/barrelShift/_0185_ ), .ZN(\EXU/ALU/barrelShift/_0203_ ) );
NOR2_X4 \EXU/ALU/barrelShift/_0727_ ( .A1(\EXU/ALU/barrelShift/_0563_ ), .A2(\EXU/ALU/barrelShift/_0547_ ), .ZN(\EXU/ALU/barrelShift/_0204_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0728_ ( .A1(\EXU/ALU/barrelShift/_0545_ ), .A2(\EXU/ALU/barrelShift/_0055_ ), .ZN(\EXU/ALU/barrelShift/_0205_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0729_ ( .A1(\EXU/ALU/barrelShift/_0544_ ), .A2(\EXU/ALU/barrelShift/_0037_ ), .ZN(\EXU/ALU/barrelShift/_0206_ ) );
AND2_X1 \EXU/ALU/barrelShift/_0730_ ( .A1(\EXU/ALU/barrelShift/_0205_ ), .A2(\EXU/ALU/barrelShift/_0206_ ), .ZN(\EXU/ALU/barrelShift/_0207_ ) );
INV_X1 \EXU/ALU/barrelShift/_0731_ ( .A(\EXU/ALU/barrelShift/_0207_ ), .ZN(\EXU/ALU/barrelShift/_0208_ ) );
OAI22_X1 \EXU/ALU/barrelShift/_0732_ ( .A1(\EXU/ALU/barrelShift/_0204_ ), .A2(\EXU/ALU/barrelShift/_0069_ ), .B1(\EXU/ALU/barrelShift/_0208_ ), .B2(\EXU/ALU/barrelShift/_0560_ ), .ZN(\EXU/ALU/barrelShift/_0209_ ) );
NOR2_X1 \EXU/ALU/barrelShift/_0733_ ( .A1(\EXU/ALU/barrelShift/_0074_ ), .A2(\EXU/ALU/barrelShift/_0163_ ), .ZN(\EXU/ALU/barrelShift/_0210_ ) );
NOR2_X2 \EXU/ALU/barrelShift/_0734_ ( .A1(\EXU/ALU/barrelShift/_0209_ ), .A2(\EXU/ALU/barrelShift/_0210_ ), .ZN(\EXU/ALU/barrelShift/_0211_ ) );
OAI22_X2 \EXU/ALU/barrelShift/_0735_ ( .A1(\EXU/ALU/barrelShift/_0211_ ), .A2(\EXU/ALU/barrelShift/_0083_ ), .B1(\EXU/ALU/barrelShift/_0562_ ), .B2(\EXU/ALU/barrelShift/_0068_ ), .ZN(\EXU/ALU/barrelShift/_0212_ ) );
OR2_X4 \EXU/ALU/barrelShift/_0736_ ( .A1(\EXU/ALU/barrelShift/_0203_ ), .A2(\EXU/ALU/barrelShift/_0212_ ), .ZN(\EXU/ALU/barrelShift/_0213_ ) );
AOI22_X1 \EXU/ALU/barrelShift/_0737_ ( .A1(\EXU/ALU/barrelShift/_0213_ ), .A2(\EXU/ALU/barrelShift/_0087_ ), .B1(\EXU/ALU/barrelShift/_0151_ ), .B2(\EXU/ALU/barrelShift/_0109_ ), .ZN(\EXU/ALU/barrelShift/_0214_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0738_ ( .A1(\EXU/ALU/barrelShift/_0202_ ), .A2(\EXU/ALU/barrelShift/_0113_ ), .A3(\EXU/ALU/barrelShift/_0214_ ), .ZN(\EXU/ALU/barrelShift/_0215_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0739_ ( .A1(\EXU/ALU/barrelShift/_0170_ ), .A2(\EXU/ALU/barrelShift/_0178_ ), .ZN(\EXU/ALU/barrelShift/_0216_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0740_ ( .A1(\EXU/ALU/barrelShift/_0201_ ), .A2(\EXU/ALU/barrelShift/_0215_ ), .A3(\EXU/ALU/barrelShift/_0216_ ), .ZN(\EXU/ALU/barrelShift/_0029_ ) );
BUF_X4 \EXU/ALU/barrelShift/_0741_ ( .A(\EXU/ALU/barrelShift/_0176_ ), .Z(\EXU/ALU/barrelShift/_0217_ ) );
AOI22_X1 \EXU/ALU/barrelShift/_0742_ ( .A1(\EXU/ALU/barrelShift/_0110_ ), .A2(\EXU/ALU/barrelShift/_0217_ ), .B1(\EXU/ALU/barrelShift/_0112_ ), .B2(\EXU/ALU/barrelShift/_0170_ ), .ZN(\EXU/ALU/barrelShift/_0218_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0743_ ( .A1(\EXU/ALU/barrelShift/_0202_ ), .A2(\EXU/ALU/barrelShift/_0197_ ), .A3(\EXU/ALU/barrelShift/_0214_ ), .ZN(\EXU/ALU/barrelShift/_0219_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0744_ ( .A1(\EXU/ALU/barrelShift/_0218_ ), .A2(\EXU/ALU/barrelShift/_0219_ ), .ZN(\EXU/ALU/barrelShift/_0028_ ) );
OAI221_X1 \EXU/ALU/barrelShift/_0745_ ( .A(\EXU/ALU/barrelShift/_0174_ ), .B1(\EXU/ALU/barrelShift/_0195_ ), .B2(\EXU/ALU/barrelShift/_0067_ ), .C1(\EXU/ALU/barrelShift/_0199_ ), .C2(\EXU/ALU/barrelShift/_0169_ ), .ZN(\EXU/ALU/barrelShift/_0220_ ) );
BUF_X4 \EXU/ALU/barrelShift/_0746_ ( .A(\EXU/ALU/barrelShift/_0086_ ), .Z(\EXU/ALU/barrelShift/_0221_ ) );
AOI221_X2 \EXU/ALU/barrelShift/_0747_ ( .A(\EXU/ALU/barrelShift/_0101_ ), .B1(\EXU/ALU/barrelShift/_0185_ ), .B2(\EXU/ALU/barrelShift/_0122_ ), .C1(\EXU/ALU/barrelShift/_0166_ ), .C2(\EXU/ALU/barrelShift/_0097_ ), .ZN(\EXU/ALU/barrelShift/_0222_ ) );
AOI221_X2 \EXU/ALU/barrelShift/_0748_ ( .A(\EXU/ALU/barrelShift/_0123_ ), .B1(\EXU/ALU/barrelShift/_0117_ ), .B2(\EXU/ALU/barrelShift/_0161_ ), .C1(\EXU/ALU/barrelShift/_0094_ ), .C2(\EXU/ALU/barrelShift/_0120_ ), .ZN(\EXU/ALU/barrelShift/_0223_ ) );
BUF_X4 \EXU/ALU/barrelShift/_0749_ ( .A(\EXU/ALU/barrelShift/_0545_ ), .Z(\EXU/ALU/barrelShift/_0224_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0750_ ( .A1(\EXU/ALU/barrelShift/_0224_ ), .A2(\EXU/ALU/barrelShift/_0051_ ), .ZN(\EXU/ALU/barrelShift/_0225_ ) );
BUF_X4 \EXU/ALU/barrelShift/_0751_ ( .A(\EXU/ALU/barrelShift/_0544_ ), .Z(\EXU/ALU/barrelShift/_0226_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0752_ ( .A1(\EXU/ALU/barrelShift/_0226_ ), .A2(\EXU/ALU/barrelShift/_0034_ ), .ZN(\EXU/ALU/barrelShift/_0227_ ) );
AND3_X1 \EXU/ALU/barrelShift/_0753_ ( .A1(\EXU/ALU/barrelShift/_0225_ ), .A2(\EXU/ALU/barrelShift/_0123_ ), .A3(\EXU/ALU/barrelShift/_0227_ ), .ZN(\EXU/ALU/barrelShift/_0228_ ) );
NOR2_X2 \EXU/ALU/barrelShift/_0754_ ( .A1(\EXU/ALU/barrelShift/_0223_ ), .A2(\EXU/ALU/barrelShift/_0228_ ), .ZN(\EXU/ALU/barrelShift/_0229_ ) );
NOR2_X1 \EXU/ALU/barrelShift/_0755_ ( .A1(\EXU/ALU/barrelShift/_0229_ ), .A2(\EXU/ALU/barrelShift/_0132_ ), .ZN(\EXU/ALU/barrelShift/_0230_ ) );
OAI21_X1 \EXU/ALU/barrelShift/_0756_ ( .A(\EXU/ALU/barrelShift/_0221_ ), .B1(\EXU/ALU/barrelShift/_0222_ ), .B2(\EXU/ALU/barrelShift/_0230_ ), .ZN(\EXU/ALU/barrelShift/_0231_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0757_ ( .A1(\EXU/ALU/barrelShift/_0220_ ), .A2(\EXU/ALU/barrelShift/_0197_ ), .A3(\EXU/ALU/barrelShift/_0231_ ), .ZN(\EXU/ALU/barrelShift/_0232_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0758_ ( .A1(\EXU/ALU/barrelShift/_0196_ ), .A2(\EXU/ALU/barrelShift/_0217_ ), .A3(\EXU/ALU/barrelShift/_0200_ ), .ZN(\EXU/ALU/barrelShift/_0233_ ) );
OAI221_X1 \EXU/ALU/barrelShift/_0759_ ( .A(\EXU/ALU/barrelShift/_0174_ ), .B1(\EXU/ALU/barrelShift/_0199_ ), .B2(\EXU/ALU/barrelShift/_0109_ ), .C1(\EXU/ALU/barrelShift/_0213_ ), .C2(\EXU/ALU/barrelShift/_0067_ ), .ZN(\EXU/ALU/barrelShift/_0234_ ) );
BUF_X4 \EXU/ALU/barrelShift/_0760_ ( .A(\EXU/ALU/barrelShift/_0112_ ), .Z(\EXU/ALU/barrelShift/_0235_ ) );
NOR2_X1 \EXU/ALU/barrelShift/_0761_ ( .A1(\EXU/ALU/barrelShift/_0104_ ), .A2(\EXU/ALU/barrelShift/_0107_ ), .ZN(\EXU/ALU/barrelShift/_0236_ ) );
AOI221_X2 \EXU/ALU/barrelShift/_0762_ ( .A(\EXU/ALU/barrelShift/_0081_ ), .B1(\EXU/ALU/barrelShift/_0236_ ), .B2(\EXU/ALU/barrelShift/_0077_ ), .C1(\EXU/ALU/barrelShift/_0185_ ), .C2(\EXU/ALU/barrelShift/_0096_ ), .ZN(\EXU/ALU/barrelShift/_0237_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0763_ ( .A1(\EXU/ALU/barrelShift/_0545_ ), .A2(\EXU/ALU/barrelShift/_0052_ ), .ZN(\EXU/ALU/barrelShift/_0238_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0764_ ( .A1(\EXU/ALU/barrelShift/_0544_ ), .A2(\EXU/ALU/barrelShift/_0035_ ), .ZN(\EXU/ALU/barrelShift/_0239_ ) );
AND2_X1 \EXU/ALU/barrelShift/_0765_ ( .A1(\EXU/ALU/barrelShift/_0238_ ), .A2(\EXU/ALU/barrelShift/_0239_ ), .ZN(\EXU/ALU/barrelShift/_0240_ ) );
INV_X1 \EXU/ALU/barrelShift/_0766_ ( .A(\EXU/ALU/barrelShift/_0240_ ), .ZN(\EXU/ALU/barrelShift/_0241_ ) );
OAI22_X2 \EXU/ALU/barrelShift/_0767_ ( .A1(\EXU/ALU/barrelShift/_0089_ ), .A2(\EXU/ALU/barrelShift/_0069_ ), .B1(\EXU/ALU/barrelShift/_0241_ ), .B2(\EXU/ALU/barrelShift/_0559_ ), .ZN(\EXU/ALU/barrelShift/_0242_ ) );
NOR2_X2 \EXU/ALU/barrelShift/_0768_ ( .A1(\EXU/ALU/barrelShift/_0093_ ), .A2(\EXU/ALU/barrelShift/_0163_ ), .ZN(\EXU/ALU/barrelShift/_0243_ ) );
NOR2_X4 \EXU/ALU/barrelShift/_0769_ ( .A1(\EXU/ALU/barrelShift/_0242_ ), .A2(\EXU/ALU/barrelShift/_0243_ ), .ZN(\EXU/ALU/barrelShift/_0244_ ) );
NOR2_X1 \EXU/ALU/barrelShift/_0770_ ( .A1(\EXU/ALU/barrelShift/_0244_ ), .A2(\EXU/ALU/barrelShift/_0132_ ), .ZN(\EXU/ALU/barrelShift/_0245_ ) );
OAI21_X1 \EXU/ALU/barrelShift/_0771_ ( .A(\EXU/ALU/barrelShift/_0221_ ), .B1(\EXU/ALU/barrelShift/_0237_ ), .B2(\EXU/ALU/barrelShift/_0245_ ), .ZN(\EXU/ALU/barrelShift/_0246_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0772_ ( .A1(\EXU/ALU/barrelShift/_0234_ ), .A2(\EXU/ALU/barrelShift/_0235_ ), .A3(\EXU/ALU/barrelShift/_0246_ ), .ZN(\EXU/ALU/barrelShift/_0247_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0773_ ( .A1(\EXU/ALU/barrelShift/_0232_ ), .A2(\EXU/ALU/barrelShift/_0233_ ), .A3(\EXU/ALU/barrelShift/_0247_ ), .ZN(\EXU/ALU/barrelShift/_0027_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0774_ ( .A1(\EXU/ALU/barrelShift/_0196_ ), .A2(\EXU/ALU/barrelShift/_0113_ ), .A3(\EXU/ALU/barrelShift/_0200_ ), .ZN(\EXU/ALU/barrelShift/_0248_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0775_ ( .A1(\EXU/ALU/barrelShift/_0234_ ), .A2(\EXU/ALU/barrelShift/_0197_ ), .A3(\EXU/ALU/barrelShift/_0246_ ), .ZN(\EXU/ALU/barrelShift/_0249_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0776_ ( .A1(\EXU/ALU/barrelShift/_0202_ ), .A2(\EXU/ALU/barrelShift/_0217_ ), .A3(\EXU/ALU/barrelShift/_0214_ ), .ZN(\EXU/ALU/barrelShift/_0250_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0777_ ( .A1(\EXU/ALU/barrelShift/_0248_ ), .A2(\EXU/ALU/barrelShift/_0249_ ), .A3(\EXU/ALU/barrelShift/_0250_ ), .ZN(\EXU/ALU/barrelShift/_0026_ ) );
OR2_X2 \EXU/ALU/barrelShift/_0778_ ( .A1(\EXU/ALU/barrelShift/_0222_ ), .A2(\EXU/ALU/barrelShift/_0230_ ), .ZN(\EXU/ALU/barrelShift/_0251_ ) );
OAI221_X1 \EXU/ALU/barrelShift/_0779_ ( .A(\EXU/ALU/barrelShift/_0174_ ), .B1(\EXU/ALU/barrelShift/_0195_ ), .B2(\EXU/ALU/barrelShift/_0198_ ), .C1(\EXU/ALU/barrelShift/_0251_ ), .C2(\EXU/ALU/barrelShift/_0067_ ), .ZN(\EXU/ALU/barrelShift/_0252_ ) );
AOI221_X1 \EXU/ALU/barrelShift/_0780_ ( .A(\EXU/ALU/barrelShift/_0101_ ), .B1(\EXU/ALU/barrelShift/_0184_ ), .B2(\EXU/ALU/barrelShift/_0185_ ), .C1(\EXU/ALU/barrelShift/_0077_ ), .C2(\EXU/ALU/barrelShift/_0193_ ), .ZN(\EXU/ALU/barrelShift/_0253_ ) );
AOI221_X1 \EXU/ALU/barrelShift/_0781_ ( .A(\EXU/ALU/barrelShift/_0558_ ), .B1(\EXU/ALU/barrelShift/_0144_ ), .B2(\EXU/ALU/barrelShift/_0161_ ), .C1(\EXU/ALU/barrelShift/_0094_ ), .C2(\EXU/ALU/barrelShift/_0147_ ), .ZN(\EXU/ALU/barrelShift/_0254_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0782_ ( .A1(\EXU/ALU/barrelShift/_0224_ ), .A2(\EXU/ALU/barrelShift/_0049_ ), .ZN(\EXU/ALU/barrelShift/_0255_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0783_ ( .A1(\EXU/ALU/barrelShift/_0226_ ), .A2(\EXU/ALU/barrelShift/_0063_ ), .ZN(\EXU/ALU/barrelShift/_0256_ ) );
AND3_X1 \EXU/ALU/barrelShift/_0784_ ( .A1(\EXU/ALU/barrelShift/_0255_ ), .A2(\EXU/ALU/barrelShift/_0123_ ), .A3(\EXU/ALU/barrelShift/_0256_ ), .ZN(\EXU/ALU/barrelShift/_0257_ ) );
NOR2_X2 \EXU/ALU/barrelShift/_0785_ ( .A1(\EXU/ALU/barrelShift/_0254_ ), .A2(\EXU/ALU/barrelShift/_0257_ ), .ZN(\EXU/ALU/barrelShift/_0258_ ) );
NOR2_X1 \EXU/ALU/barrelShift/_0786_ ( .A1(\EXU/ALU/barrelShift/_0258_ ), .A2(\EXU/ALU/barrelShift/_0132_ ), .ZN(\EXU/ALU/barrelShift/_0259_ ) );
OAI21_X1 \EXU/ALU/barrelShift/_0787_ ( .A(\EXU/ALU/barrelShift/_0221_ ), .B1(\EXU/ALU/barrelShift/_0253_ ), .B2(\EXU/ALU/barrelShift/_0259_ ), .ZN(\EXU/ALU/barrelShift/_0260_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0788_ ( .A1(\EXU/ALU/barrelShift/_0252_ ), .A2(\EXU/ALU/barrelShift/_0197_ ), .A3(\EXU/ALU/barrelShift/_0260_ ), .ZN(\EXU/ALU/barrelShift/_0261_ ) );
OR2_X4 \EXU/ALU/barrelShift/_0789_ ( .A1(\EXU/ALU/barrelShift/_0237_ ), .A2(\EXU/ALU/barrelShift/_0245_ ), .ZN(\EXU/ALU/barrelShift/_0262_ ) );
OAI221_X2 \EXU/ALU/barrelShift/_0790_ ( .A(\EXU/ALU/barrelShift/_0174_ ), .B1(\EXU/ALU/barrelShift/_0199_ ), .B2(\EXU/ALU/barrelShift/_0213_ ), .C1(\EXU/ALU/barrelShift/_0262_ ), .C2(\EXU/ALU/barrelShift/_0067_ ), .ZN(\EXU/ALU/barrelShift/_0263_ ) );
AOI221_X2 \EXU/ALU/barrelShift/_0791_ ( .A(\EXU/ALU/barrelShift/_0101_ ), .B1(\EXU/ALU/barrelShift/_0562_ ), .B2(\EXU/ALU/barrelShift/_0185_ ), .C1(\EXU/ALU/barrelShift/_0077_ ), .C2(\EXU/ALU/barrelShift/_0211_ ), .ZN(\EXU/ALU/barrelShift/_0264_ ) );
AOI221_X1 \EXU/ALU/barrelShift/_0792_ ( .A(\EXU/ALU/barrelShift/_0558_ ), .B1(\EXU/ALU/barrelShift/_0557_ ), .B2(\EXU/ALU/barrelShift/_0554_ ), .C1(\EXU/ALU/barrelShift/_0161_ ), .C2(\EXU/ALU/barrelShift/_0553_ ), .ZN(\EXU/ALU/barrelShift/_0265_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0793_ ( .A1(\EXU/ALU/barrelShift/_0224_ ), .A2(\EXU/ALU/barrelShift/_0050_ ), .ZN(\EXU/ALU/barrelShift/_0266_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0794_ ( .A1(\EXU/ALU/barrelShift/_0226_ ), .A2(\EXU/ALU/barrelShift/_0033_ ), .ZN(\EXU/ALU/barrelShift/_0267_ ) );
AND3_X1 \EXU/ALU/barrelShift/_0795_ ( .A1(\EXU/ALU/barrelShift/_0266_ ), .A2(\EXU/ALU/barrelShift/_0123_ ), .A3(\EXU/ALU/barrelShift/_0267_ ), .ZN(\EXU/ALU/barrelShift/_0268_ ) );
NOR2_X2 \EXU/ALU/barrelShift/_0796_ ( .A1(\EXU/ALU/barrelShift/_0265_ ), .A2(\EXU/ALU/barrelShift/_0268_ ), .ZN(\EXU/ALU/barrelShift/_0269_ ) );
NOR2_X1 \EXU/ALU/barrelShift/_0797_ ( .A1(\EXU/ALU/barrelShift/_0269_ ), .A2(\EXU/ALU/barrelShift/_0132_ ), .ZN(\EXU/ALU/barrelShift/_0270_ ) );
OAI21_X1 \EXU/ALU/barrelShift/_0798_ ( .A(\EXU/ALU/barrelShift/_0221_ ), .B1(\EXU/ALU/barrelShift/_0264_ ), .B2(\EXU/ALU/barrelShift/_0270_ ), .ZN(\EXU/ALU/barrelShift/_0271_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0799_ ( .A1(\EXU/ALU/barrelShift/_0263_ ), .A2(\EXU/ALU/barrelShift/_0113_ ), .A3(\EXU/ALU/barrelShift/_0271_ ), .ZN(\EXU/ALU/barrelShift/_0272_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0800_ ( .A1(\EXU/ALU/barrelShift/_0220_ ), .A2(\EXU/ALU/barrelShift/_0217_ ), .A3(\EXU/ALU/barrelShift/_0231_ ), .ZN(\EXU/ALU/barrelShift/_0273_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0801_ ( .A1(\EXU/ALU/barrelShift/_0261_ ), .A2(\EXU/ALU/barrelShift/_0272_ ), .A3(\EXU/ALU/barrelShift/_0273_ ), .ZN(\EXU/ALU/barrelShift/_0025_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0802_ ( .A1(\EXU/ALU/barrelShift/_0220_ ), .A2(\EXU/ALU/barrelShift/_0113_ ), .A3(\EXU/ALU/barrelShift/_0231_ ), .ZN(\EXU/ALU/barrelShift/_0274_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0803_ ( .A1(\EXU/ALU/barrelShift/_0263_ ), .A2(\EXU/ALU/barrelShift/_0197_ ), .A3(\EXU/ALU/barrelShift/_0271_ ), .ZN(\EXU/ALU/barrelShift/_0275_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0804_ ( .A1(\EXU/ALU/barrelShift/_0234_ ), .A2(\EXU/ALU/barrelShift/_0217_ ), .A3(\EXU/ALU/barrelShift/_0246_ ), .ZN(\EXU/ALU/barrelShift/_0276_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0805_ ( .A1(\EXU/ALU/barrelShift/_0274_ ), .A2(\EXU/ALU/barrelShift/_0275_ ), .A3(\EXU/ALU/barrelShift/_0276_ ), .ZN(\EXU/ALU/barrelShift/_0024_ ) );
OR2_X2 \EXU/ALU/barrelShift/_0806_ ( .A1(\EXU/ALU/barrelShift/_0253_ ), .A2(\EXU/ALU/barrelShift/_0259_ ), .ZN(\EXU/ALU/barrelShift/_0277_ ) );
OAI221_X2 \EXU/ALU/barrelShift/_0807_ ( .A(\EXU/ALU/barrelShift/_0174_ ), .B1(\EXU/ALU/barrelShift/_0277_ ), .B2(\EXU/ALU/barrelShift/_0067_ ), .C1(\EXU/ALU/barrelShift/_0251_ ), .C2(\EXU/ALU/barrelShift/_0199_ ), .ZN(\EXU/ALU/barrelShift/_0278_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0808_ ( .A1(\EXU/ALU/barrelShift/_0545_ ), .A2(\EXU/ALU/barrelShift/_0047_ ), .ZN(\EXU/ALU/barrelShift/_0279_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0809_ ( .A1(\EXU/ALU/barrelShift/_0544_ ), .A2(\EXU/ALU/barrelShift/_0061_ ), .ZN(\EXU/ALU/barrelShift/_0280_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0810_ ( .A1(\EXU/ALU/barrelShift/_0279_ ), .A2(\EXU/ALU/barrelShift/_0280_ ), .ZN(\EXU/ALU/barrelShift/_0281_ ) );
OAI22_X1 \EXU/ALU/barrelShift/_0811_ ( .A1(\EXU/ALU/barrelShift/_0158_ ), .A2(\EXU/ALU/barrelShift/_0069_ ), .B1(\EXU/ALU/barrelShift/_0560_ ), .B2(\EXU/ALU/barrelShift/_0281_ ), .ZN(\EXU/ALU/barrelShift/_0282_ ) );
BUF_X4 \EXU/ALU/barrelShift/_0812_ ( .A(\EXU/ALU/barrelShift/_0163_ ), .Z(\EXU/ALU/barrelShift/_0283_ ) );
NOR2_X1 \EXU/ALU/barrelShift/_0813_ ( .A1(\EXU/ALU/barrelShift/_0154_ ), .A2(\EXU/ALU/barrelShift/_0283_ ), .ZN(\EXU/ALU/barrelShift/_0284_ ) );
NOR2_X2 \EXU/ALU/barrelShift/_0814_ ( .A1(\EXU/ALU/barrelShift/_0282_ ), .A2(\EXU/ALU/barrelShift/_0284_ ), .ZN(\EXU/ALU/barrelShift/_0285_ ) );
OAI22_X2 \EXU/ALU/barrelShift/_0815_ ( .A1(\EXU/ALU/barrelShift/_0229_ ), .A2(\EXU/ALU/barrelShift/_0068_ ), .B1(\EXU/ALU/barrelShift/_0132_ ), .B2(\EXU/ALU/barrelShift/_0285_ ), .ZN(\EXU/ALU/barrelShift/_0286_ ) );
NOR3_X1 \EXU/ALU/barrelShift/_0816_ ( .A1(\EXU/ALU/barrelShift/_0160_ ), .A2(\EXU/ALU/barrelShift/_0079_ ), .A3(\EXU/ALU/barrelShift/_0164_ ), .ZN(\EXU/ALU/barrelShift/_0287_ ) );
OAI21_X1 \EXU/ALU/barrelShift/_0817_ ( .A(\EXU/ALU/barrelShift/_0221_ ), .B1(\EXU/ALU/barrelShift/_0286_ ), .B2(\EXU/ALU/barrelShift/_0287_ ), .ZN(\EXU/ALU/barrelShift/_0288_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0818_ ( .A1(\EXU/ALU/barrelShift/_0278_ ), .A2(\EXU/ALU/barrelShift/_0197_ ), .A3(\EXU/ALU/barrelShift/_0288_ ), .ZN(\EXU/ALU/barrelShift/_0289_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0819_ ( .A1(\EXU/ALU/barrelShift/_0252_ ), .A2(\EXU/ALU/barrelShift/_0217_ ), .A3(\EXU/ALU/barrelShift/_0260_ ), .ZN(\EXU/ALU/barrelShift/_0290_ ) );
OR2_X2 \EXU/ALU/barrelShift/_0820_ ( .A1(\EXU/ALU/barrelShift/_0264_ ), .A2(\EXU/ALU/barrelShift/_0270_ ), .ZN(\EXU/ALU/barrelShift/_0291_ ) );
OAI221_X2 \EXU/ALU/barrelShift/_0821_ ( .A(\EXU/ALU/barrelShift/_0174_ ), .B1(\EXU/ALU/barrelShift/_0262_ ), .B2(\EXU/ALU/barrelShift/_0198_ ), .C1(\EXU/ALU/barrelShift/_0067_ ), .C2(\EXU/ALU/barrelShift/_0291_ ), .ZN(\EXU/ALU/barrelShift/_0292_ ) );
AOI221_X1 \EXU/ALU/barrelShift/_0822_ ( .A(\EXU/ALU/barrelShift/_0081_ ), .B1(\EXU/ALU/barrelShift/_0236_ ), .B2(\EXU/ALU/barrelShift/_0078_ ), .C1(\EXU/ALU/barrelShift/_0077_ ), .C2(\EXU/ALU/barrelShift/_0244_ ), .ZN(\EXU/ALU/barrelShift/_0293_ ) );
AOI221_X1 \EXU/ALU/barrelShift/_0823_ ( .A(\EXU/ALU/barrelShift/_0558_ ), .B1(\EXU/ALU/barrelShift/_0103_ ), .B2(\EXU/ALU/barrelShift/_0161_ ), .C1(\EXU/ALU/barrelShift/_0094_ ), .C2(\EXU/ALU/barrelShift/_0106_ ), .ZN(\EXU/ALU/barrelShift/_0294_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0824_ ( .A1(\EXU/ALU/barrelShift/_0224_ ), .A2(\EXU/ALU/barrelShift/_0048_ ), .ZN(\EXU/ALU/barrelShift/_0295_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0825_ ( .A1(\EXU/ALU/barrelShift/_0226_ ), .A2(\EXU/ALU/barrelShift/_0062_ ), .ZN(\EXU/ALU/barrelShift/_0296_ ) );
AND3_X1 \EXU/ALU/barrelShift/_0826_ ( .A1(\EXU/ALU/barrelShift/_0295_ ), .A2(\EXU/ALU/barrelShift/_0123_ ), .A3(\EXU/ALU/barrelShift/_0296_ ), .ZN(\EXU/ALU/barrelShift/_0297_ ) );
NOR2_X1 \EXU/ALU/barrelShift/_0827_ ( .A1(\EXU/ALU/barrelShift/_0294_ ), .A2(\EXU/ALU/barrelShift/_0297_ ), .ZN(\EXU/ALU/barrelShift/_0298_ ) );
NOR2_X1 \EXU/ALU/barrelShift/_0828_ ( .A1(\EXU/ALU/barrelShift/_0298_ ), .A2(\EXU/ALU/barrelShift/_0132_ ), .ZN(\EXU/ALU/barrelShift/_0299_ ) );
OAI21_X1 \EXU/ALU/barrelShift/_0829_ ( .A(\EXU/ALU/barrelShift/_0221_ ), .B1(\EXU/ALU/barrelShift/_0293_ ), .B2(\EXU/ALU/barrelShift/_0299_ ), .ZN(\EXU/ALU/barrelShift/_0300_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0830_ ( .A1(\EXU/ALU/barrelShift/_0292_ ), .A2(\EXU/ALU/barrelShift/_0235_ ), .A3(\EXU/ALU/barrelShift/_0300_ ), .ZN(\EXU/ALU/barrelShift/_0301_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0831_ ( .A1(\EXU/ALU/barrelShift/_0289_ ), .A2(\EXU/ALU/barrelShift/_0290_ ), .A3(\EXU/ALU/barrelShift/_0301_ ), .ZN(\EXU/ALU/barrelShift/_0023_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0832_ ( .A1(\EXU/ALU/barrelShift/_0252_ ), .A2(\EXU/ALU/barrelShift/_0113_ ), .A3(\EXU/ALU/barrelShift/_0260_ ), .ZN(\EXU/ALU/barrelShift/_0302_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0833_ ( .A1(\EXU/ALU/barrelShift/_0292_ ), .A2(\EXU/ALU/barrelShift/_0197_ ), .A3(\EXU/ALU/barrelShift/_0300_ ), .ZN(\EXU/ALU/barrelShift/_0303_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0834_ ( .A1(\EXU/ALU/barrelShift/_0263_ ), .A2(\EXU/ALU/barrelShift/_0177_ ), .A3(\EXU/ALU/barrelShift/_0271_ ), .ZN(\EXU/ALU/barrelShift/_0304_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0835_ ( .A1(\EXU/ALU/barrelShift/_0302_ ), .A2(\EXU/ALU/barrelShift/_0303_ ), .A3(\EXU/ALU/barrelShift/_0304_ ), .ZN(\EXU/ALU/barrelShift/_0022_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0836_ ( .A1(\EXU/ALU/barrelShift/_0278_ ), .A2(\EXU/ALU/barrelShift/_0178_ ), .A3(\EXU/ALU/barrelShift/_0288_ ), .ZN(\EXU/ALU/barrelShift/_0305_ ) );
OR2_X2 \EXU/ALU/barrelShift/_0837_ ( .A1(\EXU/ALU/barrelShift/_0293_ ), .A2(\EXU/ALU/barrelShift/_0299_ ), .ZN(\EXU/ALU/barrelShift/_0306_ ) );
OAI221_X2 \EXU/ALU/barrelShift/_0838_ ( .A(\EXU/ALU/barrelShift/_0174_ ), .B1(\EXU/ALU/barrelShift/_0306_ ), .B2(\EXU/ALU/barrelShift/_0067_ ), .C1(\EXU/ALU/barrelShift/_0199_ ), .C2(\EXU/ALU/barrelShift/_0291_ ), .ZN(\EXU/ALU/barrelShift/_0307_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0839_ ( .A1(\EXU/ALU/barrelShift/_0545_ ), .A2(\EXU/ALU/barrelShift/_0046_ ), .ZN(\EXU/ALU/barrelShift/_0308_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0840_ ( .A1(\EXU/ALU/barrelShift/_0544_ ), .A2(\EXU/ALU/barrelShift/_0060_ ), .ZN(\EXU/ALU/barrelShift/_0309_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0841_ ( .A1(\EXU/ALU/barrelShift/_0308_ ), .A2(\EXU/ALU/barrelShift/_0309_ ), .ZN(\EXU/ALU/barrelShift/_0310_ ) );
OAI22_X1 \EXU/ALU/barrelShift/_0842_ ( .A1(\EXU/ALU/barrelShift/_0208_ ), .A2(\EXU/ALU/barrelShift/_0069_ ), .B1(\EXU/ALU/barrelShift/_0560_ ), .B2(\EXU/ALU/barrelShift/_0310_ ), .ZN(\EXU/ALU/barrelShift/_0311_ ) );
NOR2_X1 \EXU/ALU/barrelShift/_0843_ ( .A1(\EXU/ALU/barrelShift/_0204_ ), .A2(\EXU/ALU/barrelShift/_0283_ ), .ZN(\EXU/ALU/barrelShift/_0312_ ) );
NOR2_X2 \EXU/ALU/barrelShift/_0844_ ( .A1(\EXU/ALU/barrelShift/_0311_ ), .A2(\EXU/ALU/barrelShift/_0312_ ), .ZN(\EXU/ALU/barrelShift/_0313_ ) );
OAI22_X2 \EXU/ALU/barrelShift/_0845_ ( .A1(\EXU/ALU/barrelShift/_0269_ ), .A2(\EXU/ALU/barrelShift/_0068_ ), .B1(\EXU/ALU/barrelShift/_0313_ ), .B2(\EXU/ALU/barrelShift/_0083_ ), .ZN(\EXU/ALU/barrelShift/_0314_ ) );
BUF_X4 \EXU/ALU/barrelShift/_0846_ ( .A(\EXU/ALU/barrelShift/_0079_ ), .Z(\EXU/ALU/barrelShift/_0315_ ) );
NOR2_X1 \EXU/ALU/barrelShift/_0847_ ( .A1(\EXU/ALU/barrelShift/_0211_ ), .A2(\EXU/ALU/barrelShift/_0315_ ), .ZN(\EXU/ALU/barrelShift/_0316_ ) );
OAI21_X1 \EXU/ALU/barrelShift/_0848_ ( .A(\EXU/ALU/barrelShift/_0221_ ), .B1(\EXU/ALU/barrelShift/_0314_ ), .B2(\EXU/ALU/barrelShift/_0316_ ), .ZN(\EXU/ALU/barrelShift/_0317_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0849_ ( .A1(\EXU/ALU/barrelShift/_0307_ ), .A2(\EXU/ALU/barrelShift/_0235_ ), .A3(\EXU/ALU/barrelShift/_0317_ ), .ZN(\EXU/ALU/barrelShift/_0318_ ) );
OR3_X2 \EXU/ALU/barrelShift/_0850_ ( .A1(\EXU/ALU/barrelShift/_0286_ ), .A2(\EXU/ALU/barrelShift/_0287_ ), .A3(\EXU/ALU/barrelShift/_0067_ ), .ZN(\EXU/ALU/barrelShift/_0319_ ) );
OAI211_X2 \EXU/ALU/barrelShift/_0851_ ( .A(\EXU/ALU/barrelShift/_0174_ ), .B(\EXU/ALU/barrelShift/_0319_ ), .C1(\EXU/ALU/barrelShift/_0277_ ), .C2(\EXU/ALU/barrelShift/_0199_ ), .ZN(\EXU/ALU/barrelShift/_0320_ ) );
BUF_X4 \EXU/ALU/barrelShift/_0852_ ( .A(\EXU/ALU/barrelShift/_0115_ ), .Z(\EXU/ALU/barrelShift/_0321_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0853_ ( .A1(\EXU/ALU/barrelShift/_0224_ ), .A2(\EXU/ALU/barrelShift/_0045_ ), .ZN(\EXU/ALU/barrelShift/_0322_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0854_ ( .A1(\EXU/ALU/barrelShift/_0226_ ), .A2(\EXU/ALU/barrelShift/_0059_ ), .ZN(\EXU/ALU/barrelShift/_0323_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0855_ ( .A1(\EXU/ALU/barrelShift/_0322_ ), .A2(\EXU/ALU/barrelShift/_0323_ ), .ZN(\EXU/ALU/barrelShift/_0324_ ) );
OAI22_X1 \EXU/ALU/barrelShift/_0856_ ( .A1(\EXU/ALU/barrelShift/_0190_ ), .A2(\EXU/ALU/barrelShift/_0069_ ), .B1(\EXU/ALU/barrelShift/_0560_ ), .B2(\EXU/ALU/barrelShift/_0324_ ), .ZN(\EXU/ALU/barrelShift/_0325_ ) );
NOR2_X1 \EXU/ALU/barrelShift/_0857_ ( .A1(\EXU/ALU/barrelShift/_0135_ ), .A2(\EXU/ALU/barrelShift/_0283_ ), .ZN(\EXU/ALU/barrelShift/_0326_ ) );
NOR2_X4 \EXU/ALU/barrelShift/_0858_ ( .A1(\EXU/ALU/barrelShift/_0325_ ), .A2(\EXU/ALU/barrelShift/_0326_ ), .ZN(\EXU/ALU/barrelShift/_0327_ ) );
OAI22_X1 \EXU/ALU/barrelShift/_0859_ ( .A1(\EXU/ALU/barrelShift/_0258_ ), .A2(\EXU/ALU/barrelShift/_0068_ ), .B1(\EXU/ALU/barrelShift/_0132_ ), .B2(\EXU/ALU/barrelShift/_0327_ ), .ZN(\EXU/ALU/barrelShift/_0328_ ) );
NOR2_X1 \EXU/ALU/barrelShift/_0860_ ( .A1(\EXU/ALU/barrelShift/_0193_ ), .A2(\EXU/ALU/barrelShift/_0315_ ), .ZN(\EXU/ALU/barrelShift/_0329_ ) );
OAI21_X1 \EXU/ALU/barrelShift/_0861_ ( .A(\EXU/ALU/barrelShift/_0221_ ), .B1(\EXU/ALU/barrelShift/_0328_ ), .B2(\EXU/ALU/barrelShift/_0329_ ), .ZN(\EXU/ALU/barrelShift/_0330_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0862_ ( .A1(\EXU/ALU/barrelShift/_0320_ ), .A2(\EXU/ALU/barrelShift/_0321_ ), .A3(\EXU/ALU/barrelShift/_0330_ ), .ZN(\EXU/ALU/barrelShift/_0331_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0863_ ( .A1(\EXU/ALU/barrelShift/_0305_ ), .A2(\EXU/ALU/barrelShift/_0318_ ), .A3(\EXU/ALU/barrelShift/_0331_ ), .ZN(\EXU/ALU/barrelShift/_0021_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0864_ ( .A1(\EXU/ALU/barrelShift/_0278_ ), .A2(\EXU/ALU/barrelShift/_0113_ ), .A3(\EXU/ALU/barrelShift/_0288_ ), .ZN(\EXU/ALU/barrelShift/_0332_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0865_ ( .A1(\EXU/ALU/barrelShift/_0307_ ), .A2(\EXU/ALU/barrelShift/_0197_ ), .A3(\EXU/ALU/barrelShift/_0317_ ), .ZN(\EXU/ALU/barrelShift/_0333_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0866_ ( .A1(\EXU/ALU/barrelShift/_0292_ ), .A2(\EXU/ALU/barrelShift/_0177_ ), .A3(\EXU/ALU/barrelShift/_0300_ ), .ZN(\EXU/ALU/barrelShift/_0334_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0867_ ( .A1(\EXU/ALU/barrelShift/_0332_ ), .A2(\EXU/ALU/barrelShift/_0333_ ), .A3(\EXU/ALU/barrelShift/_0334_ ), .ZN(\EXU/ALU/barrelShift/_0020_ ) );
OR3_X2 \EXU/ALU/barrelShift/_0868_ ( .A1(\EXU/ALU/barrelShift/_0314_ ), .A2(\EXU/ALU/barrelShift/_0316_ ), .A3(\EXU/ALU/barrelShift/_0067_ ), .ZN(\EXU/ALU/barrelShift/_0335_ ) );
OAI211_X2 \EXU/ALU/barrelShift/_0869_ ( .A(\EXU/ALU/barrelShift/_0174_ ), .B(\EXU/ALU/barrelShift/_0335_ ), .C1(\EXU/ALU/barrelShift/_0306_ ), .C2(\EXU/ALU/barrelShift/_0199_ ), .ZN(\EXU/ALU/barrelShift/_0336_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0870_ ( .A1(\EXU/ALU/barrelShift/_0224_ ), .A2(\EXU/ALU/barrelShift/_0044_ ), .ZN(\EXU/ALU/barrelShift/_0337_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0871_ ( .A1(\EXU/ALU/barrelShift/_0226_ ), .A2(\EXU/ALU/barrelShift/_0058_ ), .ZN(\EXU/ALU/barrelShift/_0338_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0872_ ( .A1(\EXU/ALU/barrelShift/_0337_ ), .A2(\EXU/ALU/barrelShift/_0338_ ), .ZN(\EXU/ALU/barrelShift/_0339_ ) );
OAI22_X1 \EXU/ALU/barrelShift/_0873_ ( .A1(\EXU/ALU/barrelShift/_0241_ ), .A2(\EXU/ALU/barrelShift/_0069_ ), .B1(\EXU/ALU/barrelShift/_0560_ ), .B2(\EXU/ALU/barrelShift/_0339_ ), .ZN(\EXU/ALU/barrelShift/_0340_ ) );
NOR2_X1 \EXU/ALU/barrelShift/_0874_ ( .A1(\EXU/ALU/barrelShift/_0089_ ), .A2(\EXU/ALU/barrelShift/_0283_ ), .ZN(\EXU/ALU/barrelShift/_0341_ ) );
NOR2_X2 \EXU/ALU/barrelShift/_0875_ ( .A1(\EXU/ALU/barrelShift/_0340_ ), .A2(\EXU/ALU/barrelShift/_0341_ ), .ZN(\EXU/ALU/barrelShift/_0342_ ) );
OAI22_X1 \EXU/ALU/barrelShift/_0876_ ( .A1(\EXU/ALU/barrelShift/_0298_ ), .A2(\EXU/ALU/barrelShift/_0068_ ), .B1(\EXU/ALU/barrelShift/_0132_ ), .B2(\EXU/ALU/barrelShift/_0342_ ), .ZN(\EXU/ALU/barrelShift/_0343_ ) );
NOR2_X1 \EXU/ALU/barrelShift/_0877_ ( .A1(\EXU/ALU/barrelShift/_0244_ ), .A2(\EXU/ALU/barrelShift/_0315_ ), .ZN(\EXU/ALU/barrelShift/_0344_ ) );
OAI21_X1 \EXU/ALU/barrelShift/_0878_ ( .A(\EXU/ALU/barrelShift/_0221_ ), .B1(\EXU/ALU/barrelShift/_0343_ ), .B2(\EXU/ALU/barrelShift/_0344_ ), .ZN(\EXU/ALU/barrelShift/_0345_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0879_ ( .A1(\EXU/ALU/barrelShift/_0336_ ), .A2(\EXU/ALU/barrelShift/_0113_ ), .A3(\EXU/ALU/barrelShift/_0345_ ), .ZN(\EXU/ALU/barrelShift/_0346_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0880_ ( .A1(\EXU/ALU/barrelShift/_0320_ ), .A2(\EXU/ALU/barrelShift/_0217_ ), .A3(\EXU/ALU/barrelShift/_0330_ ), .ZN(\EXU/ALU/barrelShift/_0347_ ) );
OR2_X1 \EXU/ALU/barrelShift/_0881_ ( .A1(\EXU/ALU/barrelShift/_0328_ ), .A2(\EXU/ALU/barrelShift/_0329_ ), .ZN(\EXU/ALU/barrelShift/_0348_ ) );
NOR2_X1 \EXU/ALU/barrelShift/_0882_ ( .A1(\EXU/ALU/barrelShift/_0229_ ), .A2(\EXU/ALU/barrelShift/_0315_ ), .ZN(\EXU/ALU/barrelShift/_0349_ ) );
NOR2_X1 \EXU/ALU/barrelShift/_0883_ ( .A1(\EXU/ALU/barrelShift/_0120_ ), .A2(\EXU/ALU/barrelShift/_0283_ ), .ZN(\EXU/ALU/barrelShift/_0350_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0884_ ( .A1(\EXU/ALU/barrelShift/_0224_ ), .A2(\EXU/ALU/barrelShift/_0042_ ), .ZN(\EXU/ALU/barrelShift/_0351_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0885_ ( .A1(\EXU/ALU/barrelShift/_0226_ ), .A2(\EXU/ALU/barrelShift/_0057_ ), .ZN(\EXU/ALU/barrelShift/_0352_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0886_ ( .A1(\EXU/ALU/barrelShift/_0351_ ), .A2(\EXU/ALU/barrelShift/_0123_ ), .A3(\EXU/ALU/barrelShift/_0352_ ), .ZN(\EXU/ALU/barrelShift/_0353_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0887_ ( .A1(\EXU/ALU/barrelShift/_0225_ ), .A2(\EXU/ALU/barrelShift/_0094_ ), .A3(\EXU/ALU/barrelShift/_0227_ ), .ZN(\EXU/ALU/barrelShift/_0354_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0888_ ( .A1(\EXU/ALU/barrelShift/_0353_ ), .A2(\EXU/ALU/barrelShift/_0354_ ), .ZN(\EXU/ALU/barrelShift/_0355_ ) );
NOR2_X2 \EXU/ALU/barrelShift/_0889_ ( .A1(\EXU/ALU/barrelShift/_0350_ ), .A2(\EXU/ALU/barrelShift/_0355_ ), .ZN(\EXU/ALU/barrelShift/_0356_ ) );
OAI22_X1 \EXU/ALU/barrelShift/_0890_ ( .A1(\EXU/ALU/barrelShift/_0285_ ), .A2(\EXU/ALU/barrelShift/_0068_ ), .B1(\EXU/ALU/barrelShift/_0356_ ), .B2(\EXU/ALU/barrelShift/_0083_ ), .ZN(\EXU/ALU/barrelShift/_0357_ ) );
OR2_X2 \EXU/ALU/barrelShift/_0891_ ( .A1(\EXU/ALU/barrelShift/_0349_ ), .A2(\EXU/ALU/barrelShift/_0357_ ), .ZN(\EXU/ALU/barrelShift/_0358_ ) );
AOI22_X2 \EXU/ALU/barrelShift/_0892_ ( .A1(\EXU/ALU/barrelShift/_0348_ ), .A2(\EXU/ALU/barrelShift/_0183_ ), .B1(\EXU/ALU/barrelShift/_0358_ ), .B2(\EXU/ALU/barrelShift/_0087_ ), .ZN(\EXU/ALU/barrelShift/_0359_ ) );
BUF_X4 \EXU/ALU/barrelShift/_0893_ ( .A(\EXU/ALU/barrelShift/_0539_ ), .Z(\EXU/ALU/barrelShift/_0360_ ) );
OAI21_X1 \EXU/ALU/barrelShift/_0894_ ( .A(\EXU/ALU/barrelShift/_0360_ ), .B1(\EXU/ALU/barrelShift/_0286_ ), .B2(\EXU/ALU/barrelShift/_0287_ ), .ZN(\EXU/ALU/barrelShift/_0361_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0895_ ( .A1(\EXU/ALU/barrelShift/_0359_ ), .A2(\EXU/ALU/barrelShift/_0321_ ), .A3(\EXU/ALU/barrelShift/_0361_ ), .ZN(\EXU/ALU/barrelShift/_0362_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0896_ ( .A1(\EXU/ALU/barrelShift/_0346_ ), .A2(\EXU/ALU/barrelShift/_0347_ ), .A3(\EXU/ALU/barrelShift/_0362_ ), .ZN(\EXU/ALU/barrelShift/_0019_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0897_ ( .A1(\EXU/ALU/barrelShift/_0307_ ), .A2(\EXU/ALU/barrelShift/_0178_ ), .A3(\EXU/ALU/barrelShift/_0317_ ), .ZN(\EXU/ALU/barrelShift/_0363_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0898_ ( .A1(\EXU/ALU/barrelShift/_0320_ ), .A2(\EXU/ALU/barrelShift/_0235_ ), .A3(\EXU/ALU/barrelShift/_0330_ ), .ZN(\EXU/ALU/barrelShift/_0364_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0899_ ( .A1(\EXU/ALU/barrelShift/_0336_ ), .A2(\EXU/ALU/barrelShift/_0321_ ), .A3(\EXU/ALU/barrelShift/_0345_ ), .ZN(\EXU/ALU/barrelShift/_0365_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0900_ ( .A1(\EXU/ALU/barrelShift/_0363_ ), .A2(\EXU/ALU/barrelShift/_0364_ ), .A3(\EXU/ALU/barrelShift/_0365_ ), .ZN(\EXU/ALU/barrelShift/_0018_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0901_ ( .A1(\EXU/ALU/barrelShift/_0359_ ), .A2(\EXU/ALU/barrelShift/_0178_ ), .A3(\EXU/ALU/barrelShift/_0361_ ), .ZN(\EXU/ALU/barrelShift/_0366_ ) );
OR2_X1 \EXU/ALU/barrelShift/_0902_ ( .A1(\EXU/ALU/barrelShift/_0343_ ), .A2(\EXU/ALU/barrelShift/_0344_ ), .ZN(\EXU/ALU/barrelShift/_0367_ ) );
NOR2_X1 \EXU/ALU/barrelShift/_0903_ ( .A1(\EXU/ALU/barrelShift/_0269_ ), .A2(\EXU/ALU/barrelShift/_0315_ ), .ZN(\EXU/ALU/barrelShift/_0368_ ) );
NOR2_X1 \EXU/ALU/barrelShift/_0904_ ( .A1(\EXU/ALU/barrelShift/_0557_ ), .A2(\EXU/ALU/barrelShift/_0283_ ), .ZN(\EXU/ALU/barrelShift/_0369_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0905_ ( .A1(\EXU/ALU/barrelShift/_0224_ ), .A2(\EXU/ALU/barrelShift/_0041_ ), .ZN(\EXU/ALU/barrelShift/_0370_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0906_ ( .A1(\EXU/ALU/barrelShift/_0226_ ), .A2(\EXU/ALU/barrelShift/_0054_ ), .ZN(\EXU/ALU/barrelShift/_0371_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0907_ ( .A1(\EXU/ALU/barrelShift/_0370_ ), .A2(\EXU/ALU/barrelShift/_0123_ ), .A3(\EXU/ALU/barrelShift/_0371_ ), .ZN(\EXU/ALU/barrelShift/_0372_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0908_ ( .A1(\EXU/ALU/barrelShift/_0266_ ), .A2(\EXU/ALU/barrelShift/_0094_ ), .A3(\EXU/ALU/barrelShift/_0267_ ), .ZN(\EXU/ALU/barrelShift/_0373_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0909_ ( .A1(\EXU/ALU/barrelShift/_0372_ ), .A2(\EXU/ALU/barrelShift/_0373_ ), .ZN(\EXU/ALU/barrelShift/_0374_ ) );
NOR2_X1 \EXU/ALU/barrelShift/_0910_ ( .A1(\EXU/ALU/barrelShift/_0369_ ), .A2(\EXU/ALU/barrelShift/_0374_ ), .ZN(\EXU/ALU/barrelShift/_0375_ ) );
OAI22_X1 \EXU/ALU/barrelShift/_0911_ ( .A1(\EXU/ALU/barrelShift/_0313_ ), .A2(\EXU/ALU/barrelShift/_0068_ ), .B1(\EXU/ALU/barrelShift/_0375_ ), .B2(\EXU/ALU/barrelShift/_0083_ ), .ZN(\EXU/ALU/barrelShift/_0376_ ) );
OR2_X2 \EXU/ALU/barrelShift/_0912_ ( .A1(\EXU/ALU/barrelShift/_0368_ ), .A2(\EXU/ALU/barrelShift/_0376_ ), .ZN(\EXU/ALU/barrelShift/_0377_ ) );
AOI22_X1 \EXU/ALU/barrelShift/_0913_ ( .A1(\EXU/ALU/barrelShift/_0367_ ), .A2(\EXU/ALU/barrelShift/_0183_ ), .B1(\EXU/ALU/barrelShift/_0377_ ), .B2(\EXU/ALU/barrelShift/_0087_ ), .ZN(\EXU/ALU/barrelShift/_0378_ ) );
OAI21_X1 \EXU/ALU/barrelShift/_0914_ ( .A(\EXU/ALU/barrelShift/_0360_ ), .B1(\EXU/ALU/barrelShift/_0314_ ), .B2(\EXU/ALU/barrelShift/_0316_ ), .ZN(\EXU/ALU/barrelShift/_0379_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0915_ ( .A1(\EXU/ALU/barrelShift/_0378_ ), .A2(\EXU/ALU/barrelShift/_0235_ ), .A3(\EXU/ALU/barrelShift/_0379_ ), .ZN(\EXU/ALU/barrelShift/_0380_ ) );
NOR2_X1 \EXU/ALU/barrelShift/_0916_ ( .A1(\EXU/ALU/barrelShift/_0258_ ), .A2(\EXU/ALU/barrelShift/_0315_ ), .ZN(\EXU/ALU/barrelShift/_0381_ ) );
NOR2_X1 \EXU/ALU/barrelShift/_0917_ ( .A1(\EXU/ALU/barrelShift/_0147_ ), .A2(\EXU/ALU/barrelShift/_0283_ ), .ZN(\EXU/ALU/barrelShift/_0382_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0918_ ( .A1(\EXU/ALU/barrelShift/_0224_ ), .A2(\EXU/ALU/barrelShift/_0040_ ), .ZN(\EXU/ALU/barrelShift/_0383_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0919_ ( .A1(\EXU/ALU/barrelShift/_0226_ ), .A2(\EXU/ALU/barrelShift/_0043_ ), .ZN(\EXU/ALU/barrelShift/_0384_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0920_ ( .A1(\EXU/ALU/barrelShift/_0383_ ), .A2(\EXU/ALU/barrelShift/_0123_ ), .A3(\EXU/ALU/barrelShift/_0384_ ), .ZN(\EXU/ALU/barrelShift/_0385_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0921_ ( .A1(\EXU/ALU/barrelShift/_0255_ ), .A2(\EXU/ALU/barrelShift/_0094_ ), .A3(\EXU/ALU/barrelShift/_0256_ ), .ZN(\EXU/ALU/barrelShift/_0386_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0922_ ( .A1(\EXU/ALU/barrelShift/_0385_ ), .A2(\EXU/ALU/barrelShift/_0386_ ), .ZN(\EXU/ALU/barrelShift/_0387_ ) );
NOR2_X2 \EXU/ALU/barrelShift/_0923_ ( .A1(\EXU/ALU/barrelShift/_0382_ ), .A2(\EXU/ALU/barrelShift/_0387_ ), .ZN(\EXU/ALU/barrelShift/_0388_ ) );
OAI22_X1 \EXU/ALU/barrelShift/_0924_ ( .A1(\EXU/ALU/barrelShift/_0327_ ), .A2(\EXU/ALU/barrelShift/_0068_ ), .B1(\EXU/ALU/barrelShift/_0388_ ), .B2(\EXU/ALU/barrelShift/_0083_ ), .ZN(\EXU/ALU/barrelShift/_0389_ ) );
OR2_X1 \EXU/ALU/barrelShift/_0925_ ( .A1(\EXU/ALU/barrelShift/_0381_ ), .A2(\EXU/ALU/barrelShift/_0389_ ), .ZN(\EXU/ALU/barrelShift/_0390_ ) );
AOI22_X2 \EXU/ALU/barrelShift/_0926_ ( .A1(\EXU/ALU/barrelShift/_0183_ ), .A2(\EXU/ALU/barrelShift/_0358_ ), .B1(\EXU/ALU/barrelShift/_0390_ ), .B2(\EXU/ALU/barrelShift/_0087_ ), .ZN(\EXU/ALU/barrelShift/_0391_ ) );
OAI21_X1 \EXU/ALU/barrelShift/_0927_ ( .A(\EXU/ALU/barrelShift/_0360_ ), .B1(\EXU/ALU/barrelShift/_0328_ ), .B2(\EXU/ALU/barrelShift/_0329_ ), .ZN(\EXU/ALU/barrelShift/_0392_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0928_ ( .A1(\EXU/ALU/barrelShift/_0391_ ), .A2(\EXU/ALU/barrelShift/_0321_ ), .A3(\EXU/ALU/barrelShift/_0392_ ), .ZN(\EXU/ALU/barrelShift/_0393_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0929_ ( .A1(\EXU/ALU/barrelShift/_0366_ ), .A2(\EXU/ALU/barrelShift/_0380_ ), .A3(\EXU/ALU/barrelShift/_0393_ ), .ZN(\EXU/ALU/barrelShift/_0017_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0930_ ( .A1(\EXU/ALU/barrelShift/_0336_ ), .A2(\EXU/ALU/barrelShift/_0178_ ), .A3(\EXU/ALU/barrelShift/_0345_ ), .ZN(\EXU/ALU/barrelShift/_0394_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0931_ ( .A1(\EXU/ALU/barrelShift/_0359_ ), .A2(\EXU/ALU/barrelShift/_0235_ ), .A3(\EXU/ALU/barrelShift/_0361_ ), .ZN(\EXU/ALU/barrelShift/_0395_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0932_ ( .A1(\EXU/ALU/barrelShift/_0378_ ), .A2(\EXU/ALU/barrelShift/_0321_ ), .A3(\EXU/ALU/barrelShift/_0379_ ), .ZN(\EXU/ALU/barrelShift/_0396_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0933_ ( .A1(\EXU/ALU/barrelShift/_0394_ ), .A2(\EXU/ALU/barrelShift/_0395_ ), .A3(\EXU/ALU/barrelShift/_0396_ ), .ZN(\EXU/ALU/barrelShift/_0016_ ) );
NOR2_X1 \EXU/ALU/barrelShift/_0934_ ( .A1(\EXU/ALU/barrelShift/_0298_ ), .A2(\EXU/ALU/barrelShift/_0079_ ), .ZN(\EXU/ALU/barrelShift/_0397_ ) );
NOR2_X1 \EXU/ALU/barrelShift/_0935_ ( .A1(\EXU/ALU/barrelShift/_0106_ ), .A2(\EXU/ALU/barrelShift/_0283_ ), .ZN(\EXU/ALU/barrelShift/_0398_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0936_ ( .A1(\EXU/ALU/barrelShift/_0224_ ), .A2(\EXU/ALU/barrelShift/_0039_ ), .ZN(\EXU/ALU/barrelShift/_0399_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0937_ ( .A1(\EXU/ALU/barrelShift/_0226_ ), .A2(\EXU/ALU/barrelShift/_0032_ ), .ZN(\EXU/ALU/barrelShift/_0400_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0938_ ( .A1(\EXU/ALU/barrelShift/_0399_ ), .A2(\EXU/ALU/barrelShift/_0123_ ), .A3(\EXU/ALU/barrelShift/_0400_ ), .ZN(\EXU/ALU/barrelShift/_0401_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0939_ ( .A1(\EXU/ALU/barrelShift/_0295_ ), .A2(\EXU/ALU/barrelShift/_0094_ ), .A3(\EXU/ALU/barrelShift/_0296_ ), .ZN(\EXU/ALU/barrelShift/_0402_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0940_ ( .A1(\EXU/ALU/barrelShift/_0401_ ), .A2(\EXU/ALU/barrelShift/_0402_ ), .ZN(\EXU/ALU/barrelShift/_0403_ ) );
NOR2_X1 \EXU/ALU/barrelShift/_0941_ ( .A1(\EXU/ALU/barrelShift/_0398_ ), .A2(\EXU/ALU/barrelShift/_0403_ ), .ZN(\EXU/ALU/barrelShift/_0404_ ) );
OAI22_X1 \EXU/ALU/barrelShift/_0942_ ( .A1(\EXU/ALU/barrelShift/_0342_ ), .A2(\EXU/ALU/barrelShift/_0068_ ), .B1(\EXU/ALU/barrelShift/_0404_ ), .B2(\EXU/ALU/barrelShift/_0083_ ), .ZN(\EXU/ALU/barrelShift/_0405_ ) );
OR2_X2 \EXU/ALU/barrelShift/_0943_ ( .A1(\EXU/ALU/barrelShift/_0397_ ), .A2(\EXU/ALU/barrelShift/_0405_ ), .ZN(\EXU/ALU/barrelShift/_0406_ ) );
AOI22_X1 \EXU/ALU/barrelShift/_0944_ ( .A1(\EXU/ALU/barrelShift/_0183_ ), .A2(\EXU/ALU/barrelShift/_0377_ ), .B1(\EXU/ALU/barrelShift/_0406_ ), .B2(\EXU/ALU/barrelShift/_0087_ ), .ZN(\EXU/ALU/barrelShift/_0407_ ) );
OAI21_X1 \EXU/ALU/barrelShift/_0945_ ( .A(\EXU/ALU/barrelShift/_0360_ ), .B1(\EXU/ALU/barrelShift/_0343_ ), .B2(\EXU/ALU/barrelShift/_0344_ ), .ZN(\EXU/ALU/barrelShift/_0408_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0946_ ( .A1(\EXU/ALU/barrelShift/_0407_ ), .A2(\EXU/ALU/barrelShift/_0113_ ), .A3(\EXU/ALU/barrelShift/_0408_ ), .ZN(\EXU/ALU/barrelShift/_0409_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0947_ ( .A1(\EXU/ALU/barrelShift/_0391_ ), .A2(\EXU/ALU/barrelShift/_0217_ ), .A3(\EXU/ALU/barrelShift/_0392_ ), .ZN(\EXU/ALU/barrelShift/_0410_ ) );
NOR2_X1 \EXU/ALU/barrelShift/_0948_ ( .A1(\EXU/ALU/barrelShift/_0285_ ), .A2(\EXU/ALU/barrelShift/_0315_ ), .ZN(\EXU/ALU/barrelShift/_0411_ ) );
OR2_X1 \EXU/ALU/barrelShift/_0949_ ( .A1(\EXU/ALU/barrelShift/_0157_ ), .A2(\EXU/ALU/barrelShift/_0163_ ), .ZN(\EXU/ALU/barrelShift/_0412_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0950_ ( .A1(\EXU/ALU/barrelShift/_0281_ ), .A2(\EXU/ALU/barrelShift/_0554_ ), .ZN(\EXU/ALU/barrelShift/_0413_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0951_ ( .A1(\EXU/ALU/barrelShift/_0412_ ), .A2(\EXU/ALU/barrelShift/_0101_ ), .A3(\EXU/ALU/barrelShift/_0413_ ), .ZN(\EXU/ALU/barrelShift/_0414_ ) );
OAI21_X1 \EXU/ALU/barrelShift/_0952_ ( .A(\EXU/ALU/barrelShift/_0414_ ), .B1(\EXU/ALU/barrelShift/_0356_ ), .B2(\EXU/ALU/barrelShift/_0068_ ), .ZN(\EXU/ALU/barrelShift/_0415_ ) );
OR2_X2 \EXU/ALU/barrelShift/_0953_ ( .A1(\EXU/ALU/barrelShift/_0411_ ), .A2(\EXU/ALU/barrelShift/_0415_ ), .ZN(\EXU/ALU/barrelShift/_0416_ ) );
AOI22_X2 \EXU/ALU/barrelShift/_0954_ ( .A1(\EXU/ALU/barrelShift/_0390_ ), .A2(\EXU/ALU/barrelShift/_0183_ ), .B1(\EXU/ALU/barrelShift/_0087_ ), .B2(\EXU/ALU/barrelShift/_0416_ ), .ZN(\EXU/ALU/barrelShift/_0417_ ) );
OAI21_X1 \EXU/ALU/barrelShift/_0955_ ( .A(\EXU/ALU/barrelShift/_0360_ ), .B1(\EXU/ALU/barrelShift/_0349_ ), .B2(\EXU/ALU/barrelShift/_0357_ ), .ZN(\EXU/ALU/barrelShift/_0418_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0956_ ( .A1(\EXU/ALU/barrelShift/_0417_ ), .A2(\EXU/ALU/barrelShift/_0321_ ), .A3(\EXU/ALU/barrelShift/_0418_ ), .ZN(\EXU/ALU/barrelShift/_0419_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0957_ ( .A1(\EXU/ALU/barrelShift/_0409_ ), .A2(\EXU/ALU/barrelShift/_0410_ ), .A3(\EXU/ALU/barrelShift/_0419_ ), .ZN(\EXU/ALU/barrelShift/_0015_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0958_ ( .A1(\EXU/ALU/barrelShift/_0378_ ), .A2(\EXU/ALU/barrelShift/_0178_ ), .A3(\EXU/ALU/barrelShift/_0379_ ), .ZN(\EXU/ALU/barrelShift/_0420_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0959_ ( .A1(\EXU/ALU/barrelShift/_0407_ ), .A2(\EXU/ALU/barrelShift/_0321_ ), .A3(\EXU/ALU/barrelShift/_0408_ ), .ZN(\EXU/ALU/barrelShift/_0421_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0960_ ( .A1(\EXU/ALU/barrelShift/_0391_ ), .A2(\EXU/ALU/barrelShift/_0235_ ), .A3(\EXU/ALU/barrelShift/_0392_ ), .ZN(\EXU/ALU/barrelShift/_0422_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0961_ ( .A1(\EXU/ALU/barrelShift/_0420_ ), .A2(\EXU/ALU/barrelShift/_0421_ ), .A3(\EXU/ALU/barrelShift/_0422_ ), .ZN(\EXU/ALU/barrelShift/_0014_ ) );
NOR2_X1 \EXU/ALU/barrelShift/_0962_ ( .A1(\EXU/ALU/barrelShift/_0313_ ), .A2(\EXU/ALU/barrelShift/_0079_ ), .ZN(\EXU/ALU/barrelShift/_0423_ ) );
OR2_X1 \EXU/ALU/barrelShift/_0963_ ( .A1(\EXU/ALU/barrelShift/_0207_ ), .A2(\EXU/ALU/barrelShift/_0162_ ), .ZN(\EXU/ALU/barrelShift/_0424_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0964_ ( .A1(\EXU/ALU/barrelShift/_0310_ ), .A2(\EXU/ALU/barrelShift/_0554_ ), .ZN(\EXU/ALU/barrelShift/_0425_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0965_ ( .A1(\EXU/ALU/barrelShift/_0424_ ), .A2(\EXU/ALU/barrelShift/_0101_ ), .A3(\EXU/ALU/barrelShift/_0425_ ), .ZN(\EXU/ALU/barrelShift/_0426_ ) );
OAI21_X1 \EXU/ALU/barrelShift/_0966_ ( .A(\EXU/ALU/barrelShift/_0426_ ), .B1(\EXU/ALU/barrelShift/_0375_ ), .B2(\EXU/ALU/barrelShift/_0068_ ), .ZN(\EXU/ALU/barrelShift/_0427_ ) );
OR2_X1 \EXU/ALU/barrelShift/_0967_ ( .A1(\EXU/ALU/barrelShift/_0423_ ), .A2(\EXU/ALU/barrelShift/_0427_ ), .ZN(\EXU/ALU/barrelShift/_0428_ ) );
AOI22_X2 \EXU/ALU/barrelShift/_0968_ ( .A1(\EXU/ALU/barrelShift/_0406_ ), .A2(\EXU/ALU/barrelShift/_0151_ ), .B1(\EXU/ALU/barrelShift/_0086_ ), .B2(\EXU/ALU/barrelShift/_0428_ ), .ZN(\EXU/ALU/barrelShift/_0429_ ) );
OAI21_X1 \EXU/ALU/barrelShift/_0969_ ( .A(\EXU/ALU/barrelShift/_0360_ ), .B1(\EXU/ALU/barrelShift/_0368_ ), .B2(\EXU/ALU/barrelShift/_0376_ ), .ZN(\EXU/ALU/barrelShift/_0430_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0970_ ( .A1(\EXU/ALU/barrelShift/_0429_ ), .A2(\EXU/ALU/barrelShift/_0113_ ), .A3(\EXU/ALU/barrelShift/_0430_ ), .ZN(\EXU/ALU/barrelShift/_0431_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0971_ ( .A1(\EXU/ALU/barrelShift/_0417_ ), .A2(\EXU/ALU/barrelShift/_0217_ ), .A3(\EXU/ALU/barrelShift/_0418_ ), .ZN(\EXU/ALU/barrelShift/_0432_ ) );
NOR2_X1 \EXU/ALU/barrelShift/_0972_ ( .A1(\EXU/ALU/barrelShift/_0327_ ), .A2(\EXU/ALU/barrelShift/_0079_ ), .ZN(\EXU/ALU/barrelShift/_0433_ ) );
OR2_X1 \EXU/ALU/barrelShift/_0973_ ( .A1(\EXU/ALU/barrelShift/_0189_ ), .A2(\EXU/ALU/barrelShift/_0163_ ), .ZN(\EXU/ALU/barrelShift/_0434_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0974_ ( .A1(\EXU/ALU/barrelShift/_0324_ ), .A2(\EXU/ALU/barrelShift/_0094_ ), .ZN(\EXU/ALU/barrelShift/_0435_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0975_ ( .A1(\EXU/ALU/barrelShift/_0434_ ), .A2(\EXU/ALU/barrelShift/_0101_ ), .A3(\EXU/ALU/barrelShift/_0435_ ), .ZN(\EXU/ALU/barrelShift/_0436_ ) );
OAI21_X1 \EXU/ALU/barrelShift/_0976_ ( .A(\EXU/ALU/barrelShift/_0436_ ), .B1(\EXU/ALU/barrelShift/_0388_ ), .B2(\EXU/ALU/barrelShift/_0068_ ), .ZN(\EXU/ALU/barrelShift/_0437_ ) );
OR2_X1 \EXU/ALU/barrelShift/_0977_ ( .A1(\EXU/ALU/barrelShift/_0433_ ), .A2(\EXU/ALU/barrelShift/_0437_ ), .ZN(\EXU/ALU/barrelShift/_0438_ ) );
AOI22_X2 \EXU/ALU/barrelShift/_0978_ ( .A1(\EXU/ALU/barrelShift/_0183_ ), .A2(\EXU/ALU/barrelShift/_0416_ ), .B1(\EXU/ALU/barrelShift/_0438_ ), .B2(\EXU/ALU/barrelShift/_0086_ ), .ZN(\EXU/ALU/barrelShift/_0439_ ) );
OAI21_X1 \EXU/ALU/barrelShift/_0979_ ( .A(\EXU/ALU/barrelShift/_0360_ ), .B1(\EXU/ALU/barrelShift/_0381_ ), .B2(\EXU/ALU/barrelShift/_0389_ ), .ZN(\EXU/ALU/barrelShift/_0440_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0980_ ( .A1(\EXU/ALU/barrelShift/_0439_ ), .A2(\EXU/ALU/barrelShift/_0321_ ), .A3(\EXU/ALU/barrelShift/_0440_ ), .ZN(\EXU/ALU/barrelShift/_0441_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0981_ ( .A1(\EXU/ALU/barrelShift/_0431_ ), .A2(\EXU/ALU/barrelShift/_0432_ ), .A3(\EXU/ALU/barrelShift/_0441_ ), .ZN(\EXU/ALU/barrelShift/_0013_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0982_ ( .A1(\EXU/ALU/barrelShift/_0407_ ), .A2(\EXU/ALU/barrelShift/_0178_ ), .A3(\EXU/ALU/barrelShift/_0408_ ), .ZN(\EXU/ALU/barrelShift/_0442_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0983_ ( .A1(\EXU/ALU/barrelShift/_0417_ ), .A2(\EXU/ALU/barrelShift/_0235_ ), .A3(\EXU/ALU/barrelShift/_0418_ ), .ZN(\EXU/ALU/barrelShift/_0443_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0984_ ( .A1(\EXU/ALU/barrelShift/_0429_ ), .A2(\EXU/ALU/barrelShift/_0321_ ), .A3(\EXU/ALU/barrelShift/_0430_ ), .ZN(\EXU/ALU/barrelShift/_0444_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0985_ ( .A1(\EXU/ALU/barrelShift/_0442_ ), .A2(\EXU/ALU/barrelShift/_0443_ ), .A3(\EXU/ALU/barrelShift/_0444_ ), .ZN(\EXU/ALU/barrelShift/_0012_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0986_ ( .A1(\EXU/ALU/barrelShift/_0439_ ), .A2(\EXU/ALU/barrelShift/_0177_ ), .A3(\EXU/ALU/barrelShift/_0440_ ), .ZN(\EXU/ALU/barrelShift/_0445_ ) );
AOI21_X2 \EXU/ALU/barrelShift/_0987_ ( .A(\EXU/ALU/barrelShift/_0283_ ), .B1(\EXU/ALU/barrelShift/_0225_ ), .B2(\EXU/ALU/barrelShift/_0227_ ), .ZN(\EXU/ALU/barrelShift/_0446_ ) );
AOI21_X1 \EXU/ALU/barrelShift/_0988_ ( .A(\EXU/ALU/barrelShift/_0069_ ), .B1(\EXU/ALU/barrelShift/_0351_ ), .B2(\EXU/ALU/barrelShift/_0352_ ), .ZN(\EXU/ALU/barrelShift/_0447_ ) );
NOR3_X1 \EXU/ALU/barrelShift/_0989_ ( .A1(\EXU/ALU/barrelShift/_0446_ ), .A2(\EXU/ALU/barrelShift/_0447_ ), .A3(\EXU/ALU/barrelShift/_0083_ ), .ZN(\EXU/ALU/barrelShift/_0448_ ) );
AND2_X1 \EXU/ALU/barrelShift/_0990_ ( .A1(\EXU/ALU/barrelShift/_0412_ ), .A2(\EXU/ALU/barrelShift/_0413_ ), .ZN(\EXU/ALU/barrelShift/_0449_ ) );
AOI21_X1 \EXU/ALU/barrelShift/_0991_ ( .A(\EXU/ALU/barrelShift/_0448_ ), .B1(\EXU/ALU/barrelShift/_0449_ ), .B2(\EXU/ALU/barrelShift/_0097_ ), .ZN(\EXU/ALU/barrelShift/_0450_ ) );
OAI21_X1 \EXU/ALU/barrelShift/_0992_ ( .A(\EXU/ALU/barrelShift/_0185_ ), .B1(\EXU/ALU/barrelShift/_0350_ ), .B2(\EXU/ALU/barrelShift/_0355_ ), .ZN(\EXU/ALU/barrelShift/_0451_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0993_ ( .A1(\EXU/ALU/barrelShift/_0450_ ), .A2(\EXU/ALU/barrelShift/_0451_ ), .ZN(\EXU/ALU/barrelShift/_0452_ ) );
AOI22_X1 \EXU/ALU/barrelShift/_0994_ ( .A1(\EXU/ALU/barrelShift/_0438_ ), .A2(\EXU/ALU/barrelShift/_0151_ ), .B1(\EXU/ALU/barrelShift/_0086_ ), .B2(\EXU/ALU/barrelShift/_0452_ ), .ZN(\EXU/ALU/barrelShift/_0453_ ) );
OAI21_X1 \EXU/ALU/barrelShift/_0995_ ( .A(\EXU/ALU/barrelShift/_0539_ ), .B1(\EXU/ALU/barrelShift/_0411_ ), .B2(\EXU/ALU/barrelShift/_0415_ ), .ZN(\EXU/ALU/barrelShift/_0454_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_0996_ ( .A1(\EXU/ALU/barrelShift/_0453_ ), .A2(\EXU/ALU/barrelShift/_0115_ ), .A3(\EXU/ALU/barrelShift/_0454_ ), .ZN(\EXU/ALU/barrelShift/_0455_ ) );
NOR2_X1 \EXU/ALU/barrelShift/_0997_ ( .A1(\EXU/ALU/barrelShift/_0342_ ), .A2(\EXU/ALU/barrelShift/_0315_ ), .ZN(\EXU/ALU/barrelShift/_0456_ ) );
OR2_X1 \EXU/ALU/barrelShift/_0998_ ( .A1(\EXU/ALU/barrelShift/_0240_ ), .A2(\EXU/ALU/barrelShift/_0163_ ), .ZN(\EXU/ALU/barrelShift/_0457_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_0999_ ( .A1(\EXU/ALU/barrelShift/_0339_ ), .A2(\EXU/ALU/barrelShift/_0094_ ), .ZN(\EXU/ALU/barrelShift/_0458_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_1000_ ( .A1(\EXU/ALU/barrelShift/_0457_ ), .A2(\EXU/ALU/barrelShift/_0101_ ), .A3(\EXU/ALU/barrelShift/_0458_ ), .ZN(\EXU/ALU/barrelShift/_0459_ ) );
OAI21_X1 \EXU/ALU/barrelShift/_1001_ ( .A(\EXU/ALU/barrelShift/_0459_ ), .B1(\EXU/ALU/barrelShift/_0404_ ), .B2(\EXU/ALU/barrelShift/_0068_ ), .ZN(\EXU/ALU/barrelShift/_0460_ ) );
OAI21_X1 \EXU/ALU/barrelShift/_1002_ ( .A(\EXU/ALU/barrelShift/_0087_ ), .B1(\EXU/ALU/barrelShift/_0456_ ), .B2(\EXU/ALU/barrelShift/_0460_ ), .ZN(\EXU/ALU/barrelShift/_0461_ ) );
OAI22_X1 \EXU/ALU/barrelShift/_1003_ ( .A1(\EXU/ALU/barrelShift/_0406_ ), .A2(\EXU/ALU/barrelShift/_0198_ ), .B1(\EXU/ALU/barrelShift/_0067_ ), .B2(\EXU/ALU/barrelShift/_0428_ ), .ZN(\EXU/ALU/barrelShift/_0462_ ) );
OAI21_X2 \EXU/ALU/barrelShift/_1004_ ( .A(\EXU/ALU/barrelShift/_0461_ ), .B1(\EXU/ALU/barrelShift/_0462_ ), .B2(\EXU/ALU/barrelShift/_0221_ ), .ZN(\EXU/ALU/barrelShift/_0463_ ) );
OAI211_X2 \EXU/ALU/barrelShift/_1005_ ( .A(\EXU/ALU/barrelShift/_0445_ ), .B(\EXU/ALU/barrelShift/_0455_ ), .C1(\EXU/ALU/barrelShift/_0463_ ), .C2(\EXU/ALU/barrelShift/_0066_ ), .ZN(\EXU/ALU/barrelShift/_0011_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_1006_ ( .A1(\EXU/ALU/barrelShift/_0439_ ), .A2(\EXU/ALU/barrelShift/_0112_ ), .A3(\EXU/ALU/barrelShift/_0440_ ), .ZN(\EXU/ALU/barrelShift/_0464_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_1007_ ( .A1(\EXU/ALU/barrelShift/_0429_ ), .A2(\EXU/ALU/barrelShift/_0177_ ), .A3(\EXU/ALU/barrelShift/_0430_ ), .ZN(\EXU/ALU/barrelShift/_0465_ ) );
INV_X1 \EXU/ALU/barrelShift/_1008_ ( .A(\EXU/ALU/barrelShift/_0115_ ), .ZN(\EXU/ALU/barrelShift/_0466_ ) );
OAI211_X2 \EXU/ALU/barrelShift/_1009_ ( .A(\EXU/ALU/barrelShift/_0464_ ), .B(\EXU/ALU/barrelShift/_0465_ ), .C1(\EXU/ALU/barrelShift/_0463_ ), .C2(\EXU/ALU/barrelShift/_0466_ ), .ZN(\EXU/ALU/barrelShift/_0010_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_1010_ ( .A1(\EXU/ALU/barrelShift/_0453_ ), .A2(\EXU/ALU/barrelShift/_0178_ ), .A3(\EXU/ALU/barrelShift/_0454_ ), .ZN(\EXU/ALU/barrelShift/_0467_ ) );
OR2_X1 \EXU/ALU/barrelShift/_1011_ ( .A1(\EXU/ALU/barrelShift/_0456_ ), .A2(\EXU/ALU/barrelShift/_0460_ ), .ZN(\EXU/ALU/barrelShift/_0468_ ) );
AOI21_X1 \EXU/ALU/barrelShift/_1012_ ( .A(\EXU/ALU/barrelShift/_0283_ ), .B1(\EXU/ALU/barrelShift/_0266_ ), .B2(\EXU/ALU/barrelShift/_0267_ ), .ZN(\EXU/ALU/barrelShift/_0469_ ) );
AOI21_X1 \EXU/ALU/barrelShift/_1013_ ( .A(\EXU/ALU/barrelShift/_0069_ ), .B1(\EXU/ALU/barrelShift/_0370_ ), .B2(\EXU/ALU/barrelShift/_0371_ ), .ZN(\EXU/ALU/barrelShift/_0470_ ) );
NOR3_X1 \EXU/ALU/barrelShift/_1014_ ( .A1(\EXU/ALU/barrelShift/_0469_ ), .A2(\EXU/ALU/barrelShift/_0470_ ), .A3(\EXU/ALU/barrelShift/_0083_ ), .ZN(\EXU/ALU/barrelShift/_0471_ ) );
AND2_X1 \EXU/ALU/barrelShift/_1015_ ( .A1(\EXU/ALU/barrelShift/_0424_ ), .A2(\EXU/ALU/barrelShift/_0425_ ), .ZN(\EXU/ALU/barrelShift/_0472_ ) );
AOI21_X1 \EXU/ALU/barrelShift/_1016_ ( .A(\EXU/ALU/barrelShift/_0471_ ), .B1(\EXU/ALU/barrelShift/_0472_ ), .B2(\EXU/ALU/barrelShift/_0097_ ), .ZN(\EXU/ALU/barrelShift/_0473_ ) );
OAI21_X1 \EXU/ALU/barrelShift/_1017_ ( .A(\EXU/ALU/barrelShift/_0185_ ), .B1(\EXU/ALU/barrelShift/_0369_ ), .B2(\EXU/ALU/barrelShift/_0374_ ), .ZN(\EXU/ALU/barrelShift/_0474_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_1018_ ( .A1(\EXU/ALU/barrelShift/_0473_ ), .A2(\EXU/ALU/barrelShift/_0474_ ), .ZN(\EXU/ALU/barrelShift/_0475_ ) );
AOI22_X1 \EXU/ALU/barrelShift/_1019_ ( .A1(\EXU/ALU/barrelShift/_0468_ ), .A2(\EXU/ALU/barrelShift/_0151_ ), .B1(\EXU/ALU/barrelShift/_0086_ ), .B2(\EXU/ALU/barrelShift/_0475_ ), .ZN(\EXU/ALU/barrelShift/_0476_ ) );
OAI21_X1 \EXU/ALU/barrelShift/_1020_ ( .A(\EXU/ALU/barrelShift/_0360_ ), .B1(\EXU/ALU/barrelShift/_0423_ ), .B2(\EXU/ALU/barrelShift/_0427_ ), .ZN(\EXU/ALU/barrelShift/_0477_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_1021_ ( .A1(\EXU/ALU/barrelShift/_0476_ ), .A2(\EXU/ALU/barrelShift/_0235_ ), .A3(\EXU/ALU/barrelShift/_0477_ ), .ZN(\EXU/ALU/barrelShift/_0478_ ) );
AOI21_X1 \EXU/ALU/barrelShift/_1022_ ( .A(\EXU/ALU/barrelShift/_0163_ ), .B1(\EXU/ALU/barrelShift/_0255_ ), .B2(\EXU/ALU/barrelShift/_0256_ ), .ZN(\EXU/ALU/barrelShift/_0479_ ) );
AOI21_X1 \EXU/ALU/barrelShift/_1023_ ( .A(\EXU/ALU/barrelShift/_0069_ ), .B1(\EXU/ALU/barrelShift/_0383_ ), .B2(\EXU/ALU/barrelShift/_0384_ ), .ZN(\EXU/ALU/barrelShift/_0480_ ) );
NOR3_X1 \EXU/ALU/barrelShift/_1024_ ( .A1(\EXU/ALU/barrelShift/_0479_ ), .A2(\EXU/ALU/barrelShift/_0480_ ), .A3(\EXU/ALU/barrelShift/_0082_ ), .ZN(\EXU/ALU/barrelShift/_0481_ ) );
AND2_X1 \EXU/ALU/barrelShift/_1025_ ( .A1(\EXU/ALU/barrelShift/_0434_ ), .A2(\EXU/ALU/barrelShift/_0435_ ), .ZN(\EXU/ALU/barrelShift/_0482_ ) );
AOI21_X1 \EXU/ALU/barrelShift/_1026_ ( .A(\EXU/ALU/barrelShift/_0481_ ), .B1(\EXU/ALU/barrelShift/_0482_ ), .B2(\EXU/ALU/barrelShift/_0097_ ), .ZN(\EXU/ALU/barrelShift/_0483_ ) );
OAI21_X1 \EXU/ALU/barrelShift/_1027_ ( .A(\EXU/ALU/barrelShift/_0185_ ), .B1(\EXU/ALU/barrelShift/_0382_ ), .B2(\EXU/ALU/barrelShift/_0387_ ), .ZN(\EXU/ALU/barrelShift/_0484_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_1028_ ( .A1(\EXU/ALU/barrelShift/_0483_ ), .A2(\EXU/ALU/barrelShift/_0484_ ), .ZN(\EXU/ALU/barrelShift/_0485_ ) );
AOI22_X1 \EXU/ALU/barrelShift/_1029_ ( .A1(\EXU/ALU/barrelShift/_0183_ ), .A2(\EXU/ALU/barrelShift/_0452_ ), .B1(\EXU/ALU/barrelShift/_0485_ ), .B2(\EXU/ALU/barrelShift/_0086_ ), .ZN(\EXU/ALU/barrelShift/_0486_ ) );
OAI21_X1 \EXU/ALU/barrelShift/_1030_ ( .A(\EXU/ALU/barrelShift/_0360_ ), .B1(\EXU/ALU/barrelShift/_0433_ ), .B2(\EXU/ALU/barrelShift/_0437_ ), .ZN(\EXU/ALU/barrelShift/_0487_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_1031_ ( .A1(\EXU/ALU/barrelShift/_0486_ ), .A2(\EXU/ALU/barrelShift/_0115_ ), .A3(\EXU/ALU/barrelShift/_0487_ ), .ZN(\EXU/ALU/barrelShift/_0488_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_1032_ ( .A1(\EXU/ALU/barrelShift/_0467_ ), .A2(\EXU/ALU/barrelShift/_0478_ ), .A3(\EXU/ALU/barrelShift/_0488_ ), .ZN(\EXU/ALU/barrelShift/_0009_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_1033_ ( .A1(\EXU/ALU/barrelShift/_0476_ ), .A2(\EXU/ALU/barrelShift/_0115_ ), .A3(\EXU/ALU/barrelShift/_0477_ ), .ZN(\EXU/ALU/barrelShift/_0489_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_1034_ ( .A1(\EXU/ALU/barrelShift/_0453_ ), .A2(\EXU/ALU/barrelShift/_0112_ ), .A3(\EXU/ALU/barrelShift/_0454_ ), .ZN(\EXU/ALU/barrelShift/_0490_ ) );
OAI211_X2 \EXU/ALU/barrelShift/_1035_ ( .A(\EXU/ALU/barrelShift/_0489_ ), .B(\EXU/ALU/barrelShift/_0490_ ), .C1(\EXU/ALU/barrelShift/_0463_ ), .C2(\EXU/ALU/barrelShift/_0182_ ), .ZN(\EXU/ALU/barrelShift/_0008_ ) );
OR2_X1 \EXU/ALU/barrelShift/_1036_ ( .A1(\EXU/ALU/barrelShift/_0449_ ), .A2(\EXU/ALU/barrelShift/_0079_ ), .ZN(\EXU/ALU/barrelShift/_0491_ ) );
OAI21_X1 \EXU/ALU/barrelShift/_1037_ ( .A(\EXU/ALU/barrelShift/_0077_ ), .B1(\EXU/ALU/barrelShift/_0446_ ), .B2(\EXU/ALU/barrelShift/_0447_ ), .ZN(\EXU/ALU/barrelShift/_0492_ ) );
AND2_X1 \EXU/ALU/barrelShift/_1038_ ( .A1(\EXU/ALU/barrelShift/_0491_ ), .A2(\EXU/ALU/barrelShift/_0492_ ), .ZN(\EXU/ALU/barrelShift/_0493_ ) );
AOI22_X1 \EXU/ALU/barrelShift/_1039_ ( .A1(\EXU/ALU/barrelShift/_0493_ ), .A2(\EXU/ALU/barrelShift/_0086_ ), .B1(\EXU/ALU/barrelShift/_0151_ ), .B2(\EXU/ALU/barrelShift/_0485_ ), .ZN(\EXU/ALU/barrelShift/_0494_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_1040_ ( .A1(\EXU/ALU/barrelShift/_0452_ ), .A2(\EXU/ALU/barrelShift/_0539_ ), .ZN(\EXU/ALU/barrelShift/_0495_ ) );
AND2_X1 \EXU/ALU/barrelShift/_1041_ ( .A1(\EXU/ALU/barrelShift/_0494_ ), .A2(\EXU/ALU/barrelShift/_0495_ ), .ZN(\EXU/ALU/barrelShift/_0496_ ) );
AOI21_X1 \EXU/ALU/barrelShift/_1042_ ( .A(\EXU/ALU/barrelShift/_0163_ ), .B1(\EXU/ALU/barrelShift/_0295_ ), .B2(\EXU/ALU/barrelShift/_0296_ ), .ZN(\EXU/ALU/barrelShift/_0497_ ) );
AOI21_X1 \EXU/ALU/barrelShift/_1043_ ( .A(\EXU/ALU/barrelShift/_0069_ ), .B1(\EXU/ALU/barrelShift/_0399_ ), .B2(\EXU/ALU/barrelShift/_0400_ ), .ZN(\EXU/ALU/barrelShift/_0498_ ) );
NOR3_X1 \EXU/ALU/barrelShift/_1044_ ( .A1(\EXU/ALU/barrelShift/_0497_ ), .A2(\EXU/ALU/barrelShift/_0498_ ), .A3(\EXU/ALU/barrelShift/_0082_ ), .ZN(\EXU/ALU/barrelShift/_0499_ ) );
AND2_X1 \EXU/ALU/barrelShift/_1045_ ( .A1(\EXU/ALU/barrelShift/_0457_ ), .A2(\EXU/ALU/barrelShift/_0458_ ), .ZN(\EXU/ALU/barrelShift/_0500_ ) );
AOI21_X1 \EXU/ALU/barrelShift/_1046_ ( .A(\EXU/ALU/barrelShift/_0499_ ), .B1(\EXU/ALU/barrelShift/_0500_ ), .B2(\EXU/ALU/barrelShift/_0097_ ), .ZN(\EXU/ALU/barrelShift/_0501_ ) );
OAI21_X1 \EXU/ALU/barrelShift/_1047_ ( .A(\EXU/ALU/barrelShift/_0185_ ), .B1(\EXU/ALU/barrelShift/_0398_ ), .B2(\EXU/ALU/barrelShift/_0403_ ), .ZN(\EXU/ALU/barrelShift/_0502_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_1048_ ( .A1(\EXU/ALU/barrelShift/_0501_ ), .A2(\EXU/ALU/barrelShift/_0502_ ), .ZN(\EXU/ALU/barrelShift/_0503_ ) );
AOI22_X1 \EXU/ALU/barrelShift/_1049_ ( .A1(\EXU/ALU/barrelShift/_0151_ ), .A2(\EXU/ALU/barrelShift/_0475_ ), .B1(\EXU/ALU/barrelShift/_0503_ ), .B2(\EXU/ALU/barrelShift/_0086_ ), .ZN(\EXU/ALU/barrelShift/_0504_ ) );
OAI21_X1 \EXU/ALU/barrelShift/_1050_ ( .A(\EXU/ALU/barrelShift/_0539_ ), .B1(\EXU/ALU/barrelShift/_0456_ ), .B2(\EXU/ALU/barrelShift/_0460_ ), .ZN(\EXU/ALU/barrelShift/_0505_ ) );
AND2_X2 \EXU/ALU/barrelShift/_1051_ ( .A1(\EXU/ALU/barrelShift/_0504_ ), .A2(\EXU/ALU/barrelShift/_0505_ ), .ZN(\EXU/ALU/barrelShift/_0506_ ) );
AOI22_X1 \EXU/ALU/barrelShift/_1052_ ( .A1(\EXU/ALU/barrelShift/_0496_ ), .A2(\EXU/ALU/barrelShift/_0197_ ), .B1(\EXU/ALU/barrelShift/_0506_ ), .B2(\EXU/ALU/barrelShift/_0112_ ), .ZN(\EXU/ALU/barrelShift/_0507_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_1053_ ( .A1(\EXU/ALU/barrelShift/_0486_ ), .A2(\EXU/ALU/barrelShift/_0178_ ), .A3(\EXU/ALU/barrelShift/_0487_ ), .ZN(\EXU/ALU/barrelShift/_0508_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_1054_ ( .A1(\EXU/ALU/barrelShift/_0507_ ), .A2(\EXU/ALU/barrelShift/_0508_ ), .ZN(\EXU/ALU/barrelShift/_0007_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_1055_ ( .A1(\EXU/ALU/barrelShift/_0476_ ), .A2(\EXU/ALU/barrelShift/_0217_ ), .A3(\EXU/ALU/barrelShift/_0477_ ), .ZN(\EXU/ALU/barrelShift/_0509_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_1056_ ( .A1(\EXU/ALU/barrelShift/_0504_ ), .A2(\EXU/ALU/barrelShift/_0321_ ), .A3(\EXU/ALU/barrelShift/_0505_ ), .ZN(\EXU/ALU/barrelShift/_0510_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_1057_ ( .A1(\EXU/ALU/barrelShift/_0486_ ), .A2(\EXU/ALU/barrelShift/_0235_ ), .A3(\EXU/ALU/barrelShift/_0487_ ), .ZN(\EXU/ALU/barrelShift/_0511_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_1058_ ( .A1(\EXU/ALU/barrelShift/_0509_ ), .A2(\EXU/ALU/barrelShift/_0510_ ), .A3(\EXU/ALU/barrelShift/_0511_ ), .ZN(\EXU/ALU/barrelShift/_0006_ ) );
OAI21_X1 \EXU/ALU/barrelShift/_1059_ ( .A(\EXU/ALU/barrelShift/_0097_ ), .B1(\EXU/ALU/barrelShift/_0479_ ), .B2(\EXU/ALU/barrelShift/_0480_ ), .ZN(\EXU/ALU/barrelShift/_0512_ ) );
OAI21_X1 \EXU/ALU/barrelShift/_1060_ ( .A(\EXU/ALU/barrelShift/_0512_ ), .B1(\EXU/ALU/barrelShift/_0482_ ), .B2(\EXU/ALU/barrelShift/_0315_ ), .ZN(\EXU/ALU/barrelShift/_0513_ ) );
OAI22_X1 \EXU/ALU/barrelShift/_1061_ ( .A1(\EXU/ALU/barrelShift/_0493_ ), .A2(\EXU/ALU/barrelShift/_0067_ ), .B1(\EXU/ALU/barrelShift/_0198_ ), .B2(\EXU/ALU/barrelShift/_0485_ ), .ZN(\EXU/ALU/barrelShift/_0514_ ) );
MUX2_X2 \EXU/ALU/barrelShift/_1062_ ( .A(\EXU/ALU/barrelShift/_0513_ ), .B(\EXU/ALU/barrelShift/_0514_ ), .S(\EXU/ALU/barrelShift/_0153_ ), .Z(\EXU/ALU/barrelShift/_0515_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_1063_ ( .A1(\EXU/ALU/barrelShift/_0515_ ), .A2(\EXU/ALU/barrelShift/_0115_ ), .ZN(\EXU/ALU/barrelShift/_0516_ ) );
NAND3_X1 \EXU/ALU/barrelShift/_1064_ ( .A1(\EXU/ALU/barrelShift/_0494_ ), .A2(\EXU/ALU/barrelShift/_0177_ ), .A3(\EXU/ALU/barrelShift/_0495_ ), .ZN(\EXU/ALU/barrelShift/_0517_ ) );
OR2_X1 \EXU/ALU/barrelShift/_1065_ ( .A1(\EXU/ALU/barrelShift/_0472_ ), .A2(\EXU/ALU/barrelShift/_0079_ ), .ZN(\EXU/ALU/barrelShift/_0518_ ) );
OAI21_X1 \EXU/ALU/barrelShift/_1066_ ( .A(\EXU/ALU/barrelShift/_0077_ ), .B1(\EXU/ALU/barrelShift/_0469_ ), .B2(\EXU/ALU/barrelShift/_0470_ ), .ZN(\EXU/ALU/barrelShift/_0519_ ) );
AND2_X1 \EXU/ALU/barrelShift/_1067_ ( .A1(\EXU/ALU/barrelShift/_0518_ ), .A2(\EXU/ALU/barrelShift/_0519_ ), .ZN(\EXU/ALU/barrelShift/_0520_ ) );
AOI22_X1 \EXU/ALU/barrelShift/_1068_ ( .A1(\EXU/ALU/barrelShift/_0520_ ), .A2(\EXU/ALU/barrelShift/_0087_ ), .B1(\EXU/ALU/barrelShift/_0151_ ), .B2(\EXU/ALU/barrelShift/_0503_ ), .ZN(\EXU/ALU/barrelShift/_0521_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_1069_ ( .A1(\EXU/ALU/barrelShift/_0475_ ), .A2(\EXU/ALU/barrelShift/_0360_ ), .ZN(\EXU/ALU/barrelShift/_0522_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_1070_ ( .A1(\EXU/ALU/barrelShift/_0521_ ), .A2(\EXU/ALU/barrelShift/_0522_ ), .ZN(\EXU/ALU/barrelShift/_0523_ ) );
OAI211_X2 \EXU/ALU/barrelShift/_1071_ ( .A(\EXU/ALU/barrelShift/_0516_ ), .B(\EXU/ALU/barrelShift/_0517_ ), .C1(\EXU/ALU/barrelShift/_0066_ ), .C2(\EXU/ALU/barrelShift/_0523_ ), .ZN(\EXU/ALU/barrelShift/_0005_ ) );
AOI22_X1 \EXU/ALU/barrelShift/_1072_ ( .A1(\EXU/ALU/barrelShift/_0496_ ), .A2(\EXU/ALU/barrelShift/_0112_ ), .B1(\EXU/ALU/barrelShift/_0506_ ), .B2(\EXU/ALU/barrelShift/_0177_ ), .ZN(\EXU/ALU/barrelShift/_0524_ ) );
OAI21_X1 \EXU/ALU/barrelShift/_1073_ ( .A(\EXU/ALU/barrelShift/_0524_ ), .B1(\EXU/ALU/barrelShift/_0466_ ), .B2(\EXU/ALU/barrelShift/_0523_ ), .ZN(\EXU/ALU/barrelShift/_0004_ ) );
OAI21_X1 \EXU/ALU/barrelShift/_1074_ ( .A(\EXU/ALU/barrelShift/_0097_ ), .B1(\EXU/ALU/barrelShift/_0497_ ), .B2(\EXU/ALU/barrelShift/_0498_ ), .ZN(\EXU/ALU/barrelShift/_0525_ ) );
OAI21_X1 \EXU/ALU/barrelShift/_1075_ ( .A(\EXU/ALU/barrelShift/_0525_ ), .B1(\EXU/ALU/barrelShift/_0500_ ), .B2(\EXU/ALU/barrelShift/_0315_ ), .ZN(\EXU/ALU/barrelShift/_0526_ ) );
OAI22_X1 \EXU/ALU/barrelShift/_1076_ ( .A1(\EXU/ALU/barrelShift/_0520_ ), .A2(\EXU/ALU/barrelShift/_0067_ ), .B1(\EXU/ALU/barrelShift/_0198_ ), .B2(\EXU/ALU/barrelShift/_0503_ ), .ZN(\EXU/ALU/barrelShift/_0527_ ) );
MUX2_X1 \EXU/ALU/barrelShift/_1077_ ( .A(\EXU/ALU/barrelShift/_0526_ ), .B(\EXU/ALU/barrelShift/_0527_ ), .S(\EXU/ALU/barrelShift/_0153_ ), .Z(\EXU/ALU/barrelShift/_0528_ ) );
AOI22_X1 \EXU/ALU/barrelShift/_1078_ ( .A1(\EXU/ALU/barrelShift/_0112_ ), .A2(\EXU/ALU/barrelShift/_0528_ ), .B1(\EXU/ALU/barrelShift/_0515_ ), .B2(\EXU/ALU/barrelShift/_0177_ ), .ZN(\EXU/ALU/barrelShift/_0529_ ) );
AOI21_X1 \EXU/ALU/barrelShift/_1079_ ( .A(\EXU/ALU/barrelShift/_0198_ ), .B1(\EXU/ALU/barrelShift/_0491_ ), .B2(\EXU/ALU/barrelShift/_0492_ ), .ZN(\EXU/ALU/barrelShift/_0530_ ) );
AOI21_X1 \EXU/ALU/barrelShift/_1080_ ( .A(\EXU/ALU/barrelShift/_0530_ ), .B1(\EXU/ALU/barrelShift/_0183_ ), .B2(\EXU/ALU/barrelShift/_0513_ ), .ZN(\EXU/ALU/barrelShift/_0531_ ) );
OAI21_X1 \EXU/ALU/barrelShift/_1081_ ( .A(\EXU/ALU/barrelShift/_0529_ ), .B1(\EXU/ALU/barrelShift/_0466_ ), .B2(\EXU/ALU/barrelShift/_0531_ ), .ZN(\EXU/ALU/barrelShift/_0003_ ) );
AOI22_X1 \EXU/ALU/barrelShift/_1082_ ( .A1(\EXU/ALU/barrelShift/_0112_ ), .A2(\EXU/ALU/barrelShift/_0515_ ), .B1(\EXU/ALU/barrelShift/_0528_ ), .B2(\EXU/ALU/barrelShift/_0115_ ), .ZN(\EXU/ALU/barrelShift/_0532_ ) );
OAI21_X1 \EXU/ALU/barrelShift/_1083_ ( .A(\EXU/ALU/barrelShift/_0532_ ), .B1(\EXU/ALU/barrelShift/_0182_ ), .B2(\EXU/ALU/barrelShift/_0523_ ), .ZN(\EXU/ALU/barrelShift/_0002_ ) );
AOI21_X1 \EXU/ALU/barrelShift/_1084_ ( .A(\EXU/ALU/barrelShift/_0199_ ), .B1(\EXU/ALU/barrelShift/_0518_ ), .B2(\EXU/ALU/barrelShift/_0519_ ), .ZN(\EXU/ALU/barrelShift/_0533_ ) );
AOI21_X1 \EXU/ALU/barrelShift/_1085_ ( .A(\EXU/ALU/barrelShift/_0533_ ), .B1(\EXU/ALU/barrelShift/_0183_ ), .B2(\EXU/ALU/barrelShift/_0526_ ), .ZN(\EXU/ALU/barrelShift/_0534_ ) );
OAI22_X1 \EXU/ALU/barrelShift/_1086_ ( .A1(\EXU/ALU/barrelShift/_0534_ ), .A2(\EXU/ALU/barrelShift/_0066_ ), .B1(\EXU/ALU/barrelShift/_0531_ ), .B2(\EXU/ALU/barrelShift/_0182_ ), .ZN(\EXU/ALU/barrelShift/_0001_ ) );
NAND2_X1 \EXU/ALU/barrelShift/_1087_ ( .A1(\EXU/ALU/barrelShift/_0528_ ), .A2(\EXU/ALU/barrelShift/_0177_ ), .ZN(\EXU/ALU/barrelShift/_0535_ ) );
OAI221_X1 \EXU/ALU/barrelShift/_1088_ ( .A(\EXU/ALU/barrelShift/_0535_ ), .B1(\EXU/ALU/barrelShift/_0066_ ), .B2(\EXU/ALU/barrelShift/_0531_ ), .C1(\EXU/ALU/barrelShift/_0466_ ), .C2(\EXU/ALU/barrelShift/_0534_ ), .ZN(\EXU/ALU/barrelShift/_0000_ ) );
BUF_X1 \EXU/ALU/barrelShift/_1089_ ( .A(\EXU/ALU/barrelShift/casez_tmp_128 ), .Z(\EXU/ALU/_barrelShift_io_out [0] ) );
BUF_X1 \EXU/ALU/barrelShift/_1090_ ( .A(\EXU/ALU/barrelShift/casez_tmp_127 ), .Z(\EXU/ALU/_barrelShift_io_out [1] ) );
BUF_X1 \EXU/ALU/barrelShift/_1091_ ( .A(\EXU/ALU/barrelShift/casez_tmp_130 ), .Z(\EXU/ALU/_barrelShift_io_out [2] ) );
BUF_X1 \EXU/ALU/barrelShift/_1092_ ( .A(\EXU/ALU/barrelShift/casez_tmp_129 ), .Z(\EXU/ALU/_barrelShift_io_out [3] ) );
BUF_X1 \EXU/ALU/barrelShift/_1093_ ( .A(\EXU/ALU/barrelShift/casez_tmp_132 ), .Z(\EXU/ALU/_barrelShift_io_out [4] ) );
BUF_X1 \EXU/ALU/barrelShift/_1094_ ( .A(\EXU/ALU/barrelShift/casez_tmp_131 ), .Z(\EXU/ALU/_barrelShift_io_out [5] ) );
BUF_X1 \EXU/ALU/barrelShift/_1095_ ( .A(\EXU/ALU/barrelShift/casez_tmp_134 ), .Z(\EXU/ALU/_barrelShift_io_out [6] ) );
BUF_X1 \EXU/ALU/barrelShift/_1096_ ( .A(\EXU/ALU/barrelShift/casez_tmp_133 ), .Z(\EXU/ALU/_barrelShift_io_out [7] ) );
BUF_X1 \EXU/ALU/barrelShift/_1097_ ( .A(\EXU/ALU/barrelShift/casez_tmp_136 ), .Z(\EXU/ALU/_barrelShift_io_out [8] ) );
BUF_X1 \EXU/ALU/barrelShift/_1098_ ( .A(\EXU/ALU/barrelShift/casez_tmp_135 ), .Z(\EXU/ALU/_barrelShift_io_out [9] ) );
BUF_X1 \EXU/ALU/barrelShift/_1099_ ( .A(\EXU/ALU/barrelShift/casez_tmp_138 ), .Z(\EXU/ALU/_barrelShift_io_out [10] ) );
BUF_X1 \EXU/ALU/barrelShift/_1100_ ( .A(\EXU/ALU/barrelShift/casez_tmp_137 ), .Z(\EXU/ALU/_barrelShift_io_out [11] ) );
BUF_X1 \EXU/ALU/barrelShift/_1101_ ( .A(\EXU/ALU/barrelShift/casez_tmp_140 ), .Z(\EXU/ALU/_barrelShift_io_out [12] ) );
BUF_X1 \EXU/ALU/barrelShift/_1102_ ( .A(\EXU/ALU/barrelShift/casez_tmp_139 ), .Z(\EXU/ALU/_barrelShift_io_out [13] ) );
BUF_X1 \EXU/ALU/barrelShift/_1103_ ( .A(\EXU/ALU/barrelShift/casez_tmp_142 ), .Z(\EXU/ALU/_barrelShift_io_out [14] ) );
BUF_X1 \EXU/ALU/barrelShift/_1104_ ( .A(\EXU/ALU/barrelShift/casez_tmp_141 ), .Z(\EXU/ALU/_barrelShift_io_out [15] ) );
BUF_X1 \EXU/ALU/barrelShift/_1105_ ( .A(\EXU/ALU/barrelShift/casez_tmp_144 ), .Z(\EXU/ALU/_barrelShift_io_out [16] ) );
BUF_X1 \EXU/ALU/barrelShift/_1106_ ( .A(\EXU/ALU/barrelShift/casez_tmp_143 ), .Z(\EXU/ALU/_barrelShift_io_out [17] ) );
BUF_X1 \EXU/ALU/barrelShift/_1107_ ( .A(\EXU/ALU/barrelShift/casez_tmp_146 ), .Z(\EXU/ALU/_barrelShift_io_out [18] ) );
BUF_X1 \EXU/ALU/barrelShift/_1108_ ( .A(\EXU/ALU/barrelShift/casez_tmp_145 ), .Z(\EXU/ALU/_barrelShift_io_out [19] ) );
BUF_X1 \EXU/ALU/barrelShift/_1109_ ( .A(\EXU/ALU/barrelShift/casez_tmp_148 ), .Z(\EXU/ALU/_barrelShift_io_out [20] ) );
BUF_X1 \EXU/ALU/barrelShift/_1110_ ( .A(\EXU/ALU/barrelShift/casez_tmp_147 ), .Z(\EXU/ALU/_barrelShift_io_out [21] ) );
BUF_X1 \EXU/ALU/barrelShift/_1111_ ( .A(\EXU/ALU/barrelShift/casez_tmp_150 ), .Z(\EXU/ALU/_barrelShift_io_out [22] ) );
BUF_X1 \EXU/ALU/barrelShift/_1112_ ( .A(\EXU/ALU/barrelShift/casez_tmp_149 ), .Z(\EXU/ALU/_barrelShift_io_out [23] ) );
BUF_X1 \EXU/ALU/barrelShift/_1113_ ( .A(\EXU/ALU/barrelShift/casez_tmp_152 ), .Z(\EXU/ALU/_barrelShift_io_out [24] ) );
BUF_X1 \EXU/ALU/barrelShift/_1114_ ( .A(\EXU/ALU/barrelShift/casez_tmp_151 ), .Z(\EXU/ALU/_barrelShift_io_out [25] ) );
BUF_X1 \EXU/ALU/barrelShift/_1115_ ( .A(\EXU/ALU/barrelShift/casez_tmp_154 ), .Z(\EXU/ALU/_barrelShift_io_out [26] ) );
BUF_X1 \EXU/ALU/barrelShift/_1116_ ( .A(\EXU/ALU/barrelShift/casez_tmp_153 ), .Z(\EXU/ALU/_barrelShift_io_out [27] ) );
BUF_X1 \EXU/ALU/barrelShift/_1117_ ( .A(\EXU/ALU/barrelShift/casez_tmp_156 ), .Z(\EXU/ALU/_barrelShift_io_out [28] ) );
BUF_X1 \EXU/ALU/barrelShift/_1118_ ( .A(\EXU/ALU/barrelShift/casez_tmp_155 ), .Z(\EXU/ALU/_barrelShift_io_out [29] ) );
BUF_X1 \EXU/ALU/barrelShift/_1119_ ( .A(\EXU/ALU/barrelShift/casez_tmp_158 ), .Z(\EXU/ALU/_barrelShift_io_out [30] ) );
BUF_X1 \EXU/ALU/barrelShift/_1120_ ( .A(\EXU/ALU/barrelShift/casez_tmp_157 ), .Z(\EXU/ALU/_barrelShift_io_out [31] ) );
BUF_X1 \EXU/ALU/barrelShift/_1121_ ( .A(\EXU/casez_tmp_0 [4] ), .Z(\EXU/ALU/barrelShift/_0070_ ) );
BUF_X1 \EXU/ALU/barrelShift/_1122_ ( .A(\EXU/ALU/_aluControl_io_isLeft ), .Z(\EXU/ALU/barrelShift/_0065_ ) );
BUF_X1 \EXU/ALU/barrelShift/_1123_ ( .A(\EXU/_0006_ ), .Z(\EXU/ALU/barrelShift/_0038_ ) );
BUF_X1 \EXU/ALU/barrelShift/_1124_ ( .A(\EXU/_0024_ ), .Z(\EXU/ALU/barrelShift/_0056_ ) );
BUF_X1 \EXU/ALU/barrelShift/_1125_ ( .A(\EXU/casez_tmp_0 [3] ), .Z(\EXU/ALU/barrelShift/_0069_ ) );
BUF_X1 \EXU/ALU/barrelShift/_1126_ ( .A(\EXU/_0029_ ), .Z(\EXU/ALU/barrelShift/_0061_ ) );
BUF_X1 \EXU/ALU/barrelShift/_1127_ ( .A(\EXU/_0015_ ), .Z(\EXU/ALU/barrelShift/_0047_ ) );
BUF_X1 \EXU/ALU/barrelShift/_1128_ ( .A(\EXU/ALU/_aluControl_io_isArith ), .Z(\EXU/ALU/barrelShift/_0064_ ) );
BUF_X1 \EXU/ALU/barrelShift/_1129_ ( .A(\EXU/casez_tmp_0 [2] ), .Z(\EXU/ALU/barrelShift/_0068_ ) );
BUF_X1 \EXU/ALU/barrelShift/_1130_ ( .A(\EXU/_0025_ ), .Z(\EXU/ALU/barrelShift/_0057_ ) );
BUF_X1 \EXU/ALU/barrelShift/_1131_ ( .A(\EXU/_0010_ ), .Z(\EXU/ALU/barrelShift/_0042_ ) );
BUF_X1 \EXU/ALU/barrelShift/_1132_ ( .A(\EXU/_0002_ ), .Z(\EXU/ALU/barrelShift/_0034_ ) );
BUF_X1 \EXU/ALU/barrelShift/_1133_ ( .A(\EXU/_0019_ ), .Z(\EXU/ALU/barrelShift/_0051_ ) );
BUF_X1 \EXU/ALU/barrelShift/_1134_ ( .A(\EXU/casez_tmp_0 [1] ), .Z(\EXU/ALU/barrelShift/_0067_ ) );
BUF_X1 \EXU/ALU/barrelShift/_1135_ ( .A(\EXU/_0011_ ), .Z(\EXU/ALU/barrelShift/_0043_ ) );
BUF_X1 \EXU/ALU/barrelShift/_1136_ ( .A(\EXU/_0008_ ), .Z(\EXU/ALU/barrelShift/_0040_ ) );
BUF_X1 \EXU/ALU/barrelShift/_1137_ ( .A(\EXU/_0031_ ), .Z(\EXU/ALU/barrelShift/_0063_ ) );
BUF_X1 \EXU/ALU/barrelShift/_1138_ ( .A(\EXU/_0017_ ), .Z(\EXU/ALU/barrelShift/_0049_ ) );
BUF_X1 \EXU/ALU/barrelShift/_1139_ ( .A(\EXU/_0027_ ), .Z(\EXU/ALU/barrelShift/_0059_ ) );
BUF_X1 \EXU/ALU/barrelShift/_1140_ ( .A(\EXU/_0013_ ), .Z(\EXU/ALU/barrelShift/_0045_ ) );
BUF_X1 \EXU/ALU/barrelShift/_1141_ ( .A(\EXU/_0004_ ), .Z(\EXU/ALU/barrelShift/_0036_ ) );
BUF_X1 \EXU/ALU/barrelShift/_1142_ ( .A(\EXU/_0021_ ), .Z(\EXU/ALU/barrelShift/_0053_ ) );
BUF_X1 \EXU/ALU/barrelShift/_1143_ ( .A(\EXU/casez_tmp_0 [0] ), .Z(\EXU/ALU/barrelShift/_0066_ ) );
BUF_X1 \EXU/ALU/barrelShift/_1144_ ( .A(\EXU/_0000_ ), .Z(\EXU/ALU/barrelShift/_0032_ ) );
BUF_X1 \EXU/ALU/barrelShift/_1145_ ( .A(\EXU/_0007_ ), .Z(\EXU/ALU/barrelShift/_0039_ ) );
BUF_X1 \EXU/ALU/barrelShift/_1146_ ( .A(\EXU/_0030_ ), .Z(\EXU/ALU/barrelShift/_0062_ ) );
BUF_X1 \EXU/ALU/barrelShift/_1147_ ( .A(\EXU/_0016_ ), .Z(\EXU/ALU/barrelShift/_0048_ ) );
BUF_X1 \EXU/ALU/barrelShift/_1148_ ( .A(\EXU/_0026_ ), .Z(\EXU/ALU/barrelShift/_0058_ ) );
BUF_X1 \EXU/ALU/barrelShift/_1149_ ( .A(\EXU/_0012_ ), .Z(\EXU/ALU/barrelShift/_0044_ ) );
BUF_X1 \EXU/ALU/barrelShift/_1150_ ( .A(\EXU/_0003_ ), .Z(\EXU/ALU/barrelShift/_0035_ ) );
BUF_X1 \EXU/ALU/barrelShift/_1151_ ( .A(\EXU/_0020_ ), .Z(\EXU/ALU/barrelShift/_0052_ ) );
BUF_X1 \EXU/ALU/barrelShift/_1152_ ( .A(\EXU/_0022_ ), .Z(\EXU/ALU/barrelShift/_0054_ ) );
BUF_X1 \EXU/ALU/barrelShift/_1153_ ( .A(\EXU/_0009_ ), .Z(\EXU/ALU/barrelShift/_0041_ ) );
BUF_X1 \EXU/ALU/barrelShift/_1154_ ( .A(\EXU/_0001_ ), .Z(\EXU/ALU/barrelShift/_0033_ ) );
BUF_X1 \EXU/ALU/barrelShift/_1155_ ( .A(\EXU/_0018_ ), .Z(\EXU/ALU/barrelShift/_0050_ ) );
BUF_X1 \EXU/ALU/barrelShift/_1156_ ( .A(\EXU/_0028_ ), .Z(\EXU/ALU/barrelShift/_0060_ ) );
BUF_X1 \EXU/ALU/barrelShift/_1157_ ( .A(\EXU/_0014_ ), .Z(\EXU/ALU/barrelShift/_0046_ ) );
BUF_X1 \EXU/ALU/barrelShift/_1158_ ( .A(\EXU/_0005_ ), .Z(\EXU/ALU/barrelShift/_0037_ ) );
BUF_X1 \EXU/ALU/barrelShift/_1159_ ( .A(\EXU/_0023_ ), .Z(\EXU/ALU/barrelShift/_0055_ ) );
BUF_X1 \EXU/ALU/barrelShift/_1160_ ( .A(\EXU/ALU/barrelShift/_0031_ ), .Z(\EXU/ALU/barrelShift/casez_tmp_158 ) );
BUF_X1 \EXU/ALU/barrelShift/_1161_ ( .A(\EXU/ALU/barrelShift/_0030_ ), .Z(\EXU/ALU/barrelShift/casez_tmp_157 ) );
BUF_X1 \EXU/ALU/barrelShift/_1162_ ( .A(\EXU/ALU/barrelShift/_0029_ ), .Z(\EXU/ALU/barrelShift/casez_tmp_156 ) );
BUF_X1 \EXU/ALU/barrelShift/_1163_ ( .A(\EXU/ALU/barrelShift/_0028_ ), .Z(\EXU/ALU/barrelShift/casez_tmp_155 ) );
BUF_X1 \EXU/ALU/barrelShift/_1164_ ( .A(\EXU/ALU/barrelShift/_0027_ ), .Z(\EXU/ALU/barrelShift/casez_tmp_154 ) );
BUF_X1 \EXU/ALU/barrelShift/_1165_ ( .A(\EXU/ALU/barrelShift/_0026_ ), .Z(\EXU/ALU/barrelShift/casez_tmp_153 ) );
BUF_X1 \EXU/ALU/barrelShift/_1166_ ( .A(\EXU/ALU/barrelShift/_0025_ ), .Z(\EXU/ALU/barrelShift/casez_tmp_152 ) );
BUF_X1 \EXU/ALU/barrelShift/_1167_ ( .A(\EXU/ALU/barrelShift/_0024_ ), .Z(\EXU/ALU/barrelShift/casez_tmp_151 ) );
BUF_X1 \EXU/ALU/barrelShift/_1168_ ( .A(\EXU/ALU/barrelShift/_0023_ ), .Z(\EXU/ALU/barrelShift/casez_tmp_150 ) );
BUF_X1 \EXU/ALU/barrelShift/_1169_ ( .A(\EXU/ALU/barrelShift/_0022_ ), .Z(\EXU/ALU/barrelShift/casez_tmp_149 ) );
BUF_X1 \EXU/ALU/barrelShift/_1170_ ( .A(\EXU/ALU/barrelShift/_0021_ ), .Z(\EXU/ALU/barrelShift/casez_tmp_148 ) );
BUF_X1 \EXU/ALU/barrelShift/_1171_ ( .A(\EXU/ALU/barrelShift/_0020_ ), .Z(\EXU/ALU/barrelShift/casez_tmp_147 ) );
BUF_X1 \EXU/ALU/barrelShift/_1172_ ( .A(\EXU/ALU/barrelShift/_0019_ ), .Z(\EXU/ALU/barrelShift/casez_tmp_146 ) );
BUF_X1 \EXU/ALU/barrelShift/_1173_ ( .A(\EXU/ALU/barrelShift/_0018_ ), .Z(\EXU/ALU/barrelShift/casez_tmp_145 ) );
BUF_X1 \EXU/ALU/barrelShift/_1174_ ( .A(\EXU/ALU/barrelShift/_0017_ ), .Z(\EXU/ALU/barrelShift/casez_tmp_144 ) );
BUF_X1 \EXU/ALU/barrelShift/_1175_ ( .A(\EXU/ALU/barrelShift/_0016_ ), .Z(\EXU/ALU/barrelShift/casez_tmp_143 ) );
BUF_X1 \EXU/ALU/barrelShift/_1176_ ( .A(\EXU/ALU/barrelShift/_0015_ ), .Z(\EXU/ALU/barrelShift/casez_tmp_142 ) );
BUF_X1 \EXU/ALU/barrelShift/_1177_ ( .A(\EXU/ALU/barrelShift/_0014_ ), .Z(\EXU/ALU/barrelShift/casez_tmp_141 ) );
BUF_X1 \EXU/ALU/barrelShift/_1178_ ( .A(\EXU/ALU/barrelShift/_0013_ ), .Z(\EXU/ALU/barrelShift/casez_tmp_140 ) );
BUF_X1 \EXU/ALU/barrelShift/_1179_ ( .A(\EXU/ALU/barrelShift/_0012_ ), .Z(\EXU/ALU/barrelShift/casez_tmp_139 ) );
BUF_X1 \EXU/ALU/barrelShift/_1180_ ( .A(\EXU/ALU/barrelShift/_0011_ ), .Z(\EXU/ALU/barrelShift/casez_tmp_138 ) );
BUF_X1 \EXU/ALU/barrelShift/_1181_ ( .A(\EXU/ALU/barrelShift/_0010_ ), .Z(\EXU/ALU/barrelShift/casez_tmp_137 ) );
BUF_X1 \EXU/ALU/barrelShift/_1182_ ( .A(\EXU/ALU/barrelShift/_0009_ ), .Z(\EXU/ALU/barrelShift/casez_tmp_136 ) );
BUF_X1 \EXU/ALU/barrelShift/_1183_ ( .A(\EXU/ALU/barrelShift/_0008_ ), .Z(\EXU/ALU/barrelShift/casez_tmp_135 ) );
BUF_X1 \EXU/ALU/barrelShift/_1184_ ( .A(\EXU/ALU/barrelShift/_0007_ ), .Z(\EXU/ALU/barrelShift/casez_tmp_134 ) );
BUF_X1 \EXU/ALU/barrelShift/_1185_ ( .A(\EXU/ALU/barrelShift/_0006_ ), .Z(\EXU/ALU/barrelShift/casez_tmp_133 ) );
BUF_X1 \EXU/ALU/barrelShift/_1186_ ( .A(\EXU/ALU/barrelShift/_0005_ ), .Z(\EXU/ALU/barrelShift/casez_tmp_132 ) );
BUF_X1 \EXU/ALU/barrelShift/_1187_ ( .A(\EXU/ALU/barrelShift/_0004_ ), .Z(\EXU/ALU/barrelShift/casez_tmp_131 ) );
BUF_X1 \EXU/ALU/barrelShift/_1188_ ( .A(\EXU/ALU/barrelShift/_0003_ ), .Z(\EXU/ALU/barrelShift/casez_tmp_130 ) );
BUF_X1 \EXU/ALU/barrelShift/_1189_ ( .A(\EXU/ALU/barrelShift/_0002_ ), .Z(\EXU/ALU/barrelShift/casez_tmp_129 ) );
BUF_X1 \EXU/ALU/barrelShift/_1190_ ( .A(\EXU/ALU/barrelShift/_0001_ ), .Z(\EXU/ALU/barrelShift/casez_tmp_128 ) );
BUF_X1 \EXU/ALU/barrelShift/_1191_ ( .A(\EXU/ALU/barrelShift/_0000_ ), .Z(\EXU/ALU/barrelShift/casez_tmp_127 ) );
INV_X32 \EXU/BrCond/_17_ ( .A(\EXU/BrCond/_03_ ), .ZN(\EXU/BrCond/_16_ ) );
OR3_X2 \EXU/BrCond/_18_ ( .A1(\EXU/BrCond/_16_ ), .A2(\EXU/BrCond/_04_ ), .A3(\EXU/BrCond/_02_ ), .ZN(\EXU/BrCond/_01_ ) );
NAND3_X1 \EXU/BrCond/_19_ ( .A1(\EXU/BrCond/_16_ ), .A2(\EXU/BrCond/_04_ ), .A3(\EXU/BrCond/_02_ ), .ZN(\EXU/BrCond/_07_ ) );
NOR2_X1 \EXU/BrCond/_20_ ( .A1(\EXU/BrCond/_07_ ), .A2(\EXU/BrCond/_06_ ), .ZN(\EXU/BrCond/_08_ ) );
INV_X32 \EXU/BrCond/_21_ ( .A(\EXU/BrCond/_02_ ), .ZN(\EXU/BrCond/_09_ ) );
AND4_X4 \EXU/BrCond/_22_ ( .A1(\EXU/BrCond/_04_ ), .A2(\EXU/BrCond/_09_ ), .A3(\EXU/BrCond/_03_ ), .A4(\EXU/BrCond/_05_ ), .ZN(\EXU/BrCond/_10_ ) );
NAND3_X2 \EXU/BrCond/_23_ ( .A1(\EXU/BrCond/_04_ ), .A2(\EXU/BrCond/_02_ ), .A3(\EXU/BrCond/_03_ ), .ZN(\EXU/BrCond/_11_ ) );
NOR2_X1 \EXU/BrCond/_24_ ( .A1(\EXU/BrCond/_11_ ), .A2(\EXU/BrCond/_05_ ), .ZN(\EXU/BrCond/_12_ ) );
NOR3_X2 \EXU/BrCond/_25_ ( .A1(\EXU/BrCond/_08_ ), .A2(\EXU/BrCond/_10_ ), .A3(\EXU/BrCond/_12_ ), .ZN(\EXU/BrCond/_13_ ) );
NAND4_X1 \EXU/BrCond/_26_ ( .A1(\EXU/BrCond/_09_ ), .A2(\EXU/BrCond/_16_ ), .A3(\EXU/BrCond/_04_ ), .A4(\EXU/BrCond/_06_ ), .ZN(\EXU/BrCond/_14_ ) );
OR3_X4 \EXU/BrCond/_27_ ( .A1(\EXU/BrCond/_09_ ), .A2(\EXU/BrCond/_04_ ), .A3(\EXU/BrCond/_03_ ), .ZN(\EXU/BrCond/_15_ ) );
NAND4_X1 \EXU/BrCond/_28_ ( .A1(\EXU/BrCond/_13_ ), .A2(\EXU/BrCond/_01_ ), .A3(\EXU/BrCond/_14_ ), .A4(\EXU/BrCond/_15_ ), .ZN(\EXU/BrCond/_00_ ) );
BUF_X1 \EXU/BrCond/_29_ ( .A(\EXU/in_control_brType [2] ), .Z(\EXU/BrCond/_04_ ) );
BUF_X1 \EXU/BrCond/_30_ ( .A(\EXU/in_control_brType [0] ), .Z(\EXU/BrCond/_02_ ) );
BUF_X1 \EXU/BrCond/_31_ ( .A(\EXU/in_control_brType [1] ), .Z(\EXU/BrCond/_03_ ) );
BUF_X1 \EXU/BrCond/_32_ ( .A(\EXU/BrCond/_01_ ), .Z(\EXU/_BrCond_io_PCBSrc ) );
BUF_X1 \EXU/BrCond/_33_ ( .A(\EXU/_ALU_io_zero ), .Z(\EXU/BrCond/_06_ ) );
BUF_X1 \EXU/BrCond/_34_ ( .A(\EXU/_ALU_io_less ), .Z(\EXU/BrCond/_05_ ) );
BUF_X1 \EXU/BrCond/_35_ ( .A(\EXU/BrCond/_00_ ), .Z(\EXU/_BrCond_io_PCASrc ) );
NOR2_X1 \EXU/CSRControl/_1634_ ( .A1(fanout_net_18 ), .A2(fanout_net_17 ), .ZN(\EXU/CSRControl/_0795_ ) );
INV_X32 \EXU/CSRControl/_1635_ ( .A(\EXU/CSRControl/_0274_ ), .ZN(\EXU/CSRControl/_0796_ ) );
AND2_X2 \EXU/CSRControl/_1636_ ( .A1(\EXU/CSRControl/_0795_ ), .A2(\EXU/CSRControl/_0796_ ), .ZN(\EXU/CSRControl/_0797_ ) );
BUF_X4 \EXU/CSRControl/_1637_ ( .A(\EXU/CSRControl/_0797_ ), .Z(\EXU/CSRControl/_0798_ ) );
BUF_X4 \EXU/CSRControl/_1638_ ( .A(\EXU/CSRControl/_0796_ ), .Z(\EXU/CSRControl/_0799_ ) );
BUF_X4 \EXU/CSRControl/_1639_ ( .A(\EXU/CSRControl/_0799_ ), .Z(\EXU/CSRControl/_0800_ ) );
BUF_X4 \EXU/CSRControl/_1640_ ( .A(\EXU/CSRControl/_0800_ ), .Z(\EXU/CSRControl/_0801_ ) );
NOR4_X1 \EXU/CSRControl/_1641_ ( .A1(\EXU/CSRControl/_0801_ ), .A2(fanout_net_18 ), .A3(fanout_net_17 ), .A4(\EXU/CSRControl/_0164_ ), .ZN(\EXU/CSRControl/_0802_ ) );
NOR2_X4 \EXU/CSRControl/_1642_ ( .A1(\EXU/CSRControl/_0796_ ), .A2(fanout_net_18 ), .ZN(\EXU/CSRControl/_0803_ ) );
AND2_X2 \EXU/CSRControl/_1643_ ( .A1(\EXU/CSRControl/_0803_ ), .A2(fanout_net_17 ), .ZN(\EXU/CSRControl/_0804_ ) );
BUF_X4 \EXU/CSRControl/_1644_ ( .A(\EXU/CSRControl/_0804_ ), .Z(\EXU/CSRControl/_0805_ ) );
INV_X1 \EXU/CSRControl/_1645_ ( .A(\EXU/CSRControl/_0265_ ), .ZN(\EXU/CSRControl/_0806_ ) );
NOR2_X4 \EXU/CSRControl/_1646_ ( .A1(\EXU/CSRControl/_0267_ ), .A2(\EXU/CSRControl/_0266_ ), .ZN(\EXU/CSRControl/_0807_ ) );
NOR2_X4 \EXU/CSRControl/_1647_ ( .A1(\EXU/CSRControl/_0269_ ), .A2(\EXU/CSRControl/_0268_ ), .ZN(\EXU/CSRControl/_0808_ ) );
AND2_X4 \EXU/CSRControl/_1648_ ( .A1(\EXU/CSRControl/_0807_ ), .A2(\EXU/CSRControl/_0808_ ), .ZN(\EXU/CSRControl/_0809_ ) );
INV_X16 \EXU/CSRControl/_1649_ ( .A(\EXU/CSRControl/_0260_ ), .ZN(\EXU/CSRControl/_0810_ ) );
NOR2_X4 \EXU/CSRControl/_1650_ ( .A1(\EXU/CSRControl/_0810_ ), .A2(\EXU/CSRControl/_0263_ ), .ZN(\EXU/CSRControl/_0811_ ) );
AND4_X4 \EXU/CSRControl/_1651_ ( .A1(\EXU/CSRControl/_0806_ ), .A2(\EXU/CSRControl/_0809_ ), .A3(\EXU/CSRControl/_0264_ ), .A4(\EXU/CSRControl/_0811_ ), .ZN(\EXU/CSRControl/_0812_ ) );
BUF_X4 \EXU/CSRControl/_1652_ ( .A(\EXU/CSRControl/_0812_ ), .Z(\EXU/CSRControl/_0813_ ) );
AND2_X4 \EXU/CSRControl/_1653_ ( .A1(\EXU/CSRControl/_0271_ ), .A2(\EXU/CSRControl/_0270_ ), .ZN(\EXU/CSRControl/_0814_ ) );
BUF_X4 \EXU/CSRControl/_1654_ ( .A(\EXU/CSRControl/_0814_ ), .Z(\EXU/CSRControl/_0815_ ) );
BUF_X4 \EXU/CSRControl/_1655_ ( .A(\EXU/CSRControl/_0815_ ), .Z(\EXU/CSRControl/_0816_ ) );
NAND3_X1 \EXU/CSRControl/_1656_ ( .A1(\EXU/CSRControl/_0813_ ), .A2(\EXU/CSRControl/_0164_ ), .A3(\EXU/CSRControl/_0816_ ), .ZN(\EXU/CSRControl/_0817_ ) );
NOR2_X4 \EXU/CSRControl/_1657_ ( .A1(\EXU/CSRControl/_0265_ ), .A2(\EXU/CSRControl/_0264_ ), .ZN(\EXU/CSRControl/_0818_ ) );
NOR2_X2 \EXU/CSRControl/_1658_ ( .A1(\EXU/CSRControl/_0263_ ), .A2(\EXU/CSRControl/_0260_ ), .ZN(\EXU/CSRControl/_0819_ ) );
AND4_X2 \EXU/CSRControl/_1659_ ( .A1(\EXU/CSRControl/_0807_ ), .A2(\EXU/CSRControl/_0818_ ), .A3(\EXU/CSRControl/_0808_ ), .A4(\EXU/CSRControl/_0819_ ), .ZN(\EXU/CSRControl/_0820_ ) );
BUF_X4 \EXU/CSRControl/_1660_ ( .A(\EXU/CSRControl/_0820_ ), .Z(\EXU/CSRControl/_0821_ ) );
BUF_X2 \EXU/CSRControl/_1661_ ( .A(\EXU/CSRControl/_0815_ ), .Z(\EXU/CSRControl/_0822_ ) );
NAND3_X1 \EXU/CSRControl/_1662_ ( .A1(\EXU/CSRControl/_0821_ ), .A2(\EXU/CSRControl/_0228_ ), .A3(\EXU/CSRControl/_0822_ ), .ZN(\EXU/CSRControl/_0823_ ) );
NAND2_X4 \EXU/CSRControl/_1663_ ( .A1(\EXU/CSRControl/_0807_ ), .A2(\EXU/CSRControl/_0268_ ), .ZN(\EXU/CSRControl/_0824_ ) );
NOR2_X4 \EXU/CSRControl/_1664_ ( .A1(\EXU/CSRControl/_0824_ ), .A2(\EXU/CSRControl/_0269_ ), .ZN(\EXU/CSRControl/_0825_ ) );
BUF_X8 \EXU/CSRControl/_1665_ ( .A(\EXU/CSRControl/_0825_ ), .Z(\EXU/CSRControl/_0826_ ) );
BUF_X4 \EXU/CSRControl/_1666_ ( .A(\EXU/CSRControl/_0826_ ), .Z(\EXU/CSRControl/_0827_ ) );
AND2_X2 \EXU/CSRControl/_1667_ ( .A1(\EXU/CSRControl/_0811_ ), .A2(\EXU/CSRControl/_0818_ ), .ZN(\EXU/CSRControl/_0828_ ) );
BUF_X4 \EXU/CSRControl/_1668_ ( .A(\EXU/CSRControl/_0828_ ), .Z(\EXU/CSRControl/_0829_ ) );
BUF_X4 \EXU/CSRControl/_1669_ ( .A(\EXU/CSRControl/_0815_ ), .Z(\EXU/CSRControl/_0830_ ) );
NAND4_X1 \EXU/CSRControl/_1670_ ( .A1(\EXU/CSRControl/_0827_ ), .A2(\EXU/CSRControl/_0829_ ), .A3(\EXU/CSRControl/_0196_ ), .A4(\EXU/CSRControl/_0830_ ), .ZN(\EXU/CSRControl/_0831_ ) );
AND3_X1 \EXU/CSRControl/_1671_ ( .A1(\EXU/CSRControl/_0817_ ), .A2(\EXU/CSRControl/_0823_ ), .A3(\EXU/CSRControl/_0831_ ), .ZN(\EXU/CSRControl/_0832_ ) );
AND4_X2 \EXU/CSRControl/_1672_ ( .A1(\EXU/CSRControl/_0263_ ), .A2(\EXU/CSRControl/_0825_ ), .A3(\EXU/CSRControl/_0810_ ), .A4(\EXU/CSRControl/_0818_ ), .ZN(\EXU/CSRControl/_0833_ ) );
BUF_X4 \EXU/CSRControl/_1673_ ( .A(\EXU/CSRControl/_0833_ ), .Z(\EXU/CSRControl/_0834_ ) );
BUF_X4 \EXU/CSRControl/_1674_ ( .A(\EXU/CSRControl/_0816_ ), .Z(\EXU/CSRControl/_0835_ ) );
NAND3_X1 \EXU/CSRControl/_1675_ ( .A1(\EXU/CSRControl/_0834_ ), .A2(\EXU/CSRControl/_0132_ ), .A3(\EXU/CSRControl/_0835_ ), .ZN(\EXU/CSRControl/_0836_ ) );
AOI21_X1 \EXU/CSRControl/_1676_ ( .A(\EXU/CSRControl/_0805_ ), .B1(\EXU/CSRControl/_0832_ ), .B2(\EXU/CSRControl/_0836_ ), .ZN(\EXU/CSRControl/_0837_ ) );
BUF_X4 \EXU/CSRControl/_1677_ ( .A(\EXU/CSRControl/_0805_ ), .Z(\EXU/CSRControl/_0838_ ) );
AOI21_X1 \EXU/CSRControl/_1678_ ( .A(\EXU/CSRControl/_0837_ ), .B1(\EXU/CSRControl/_0196_ ), .B2(\EXU/CSRControl/_0838_ ), .ZN(\EXU/CSRControl/_0839_ ) );
AND2_X1 \EXU/CSRControl/_1679_ ( .A1(\EXU/CSRControl/_0795_ ), .A2(\EXU/CSRControl/_0274_ ), .ZN(\EXU/CSRControl/_0840_ ) );
BUF_X4 \EXU/CSRControl/_1680_ ( .A(\EXU/CSRControl/_0840_ ), .Z(\EXU/CSRControl/_0841_ ) );
INV_X1 \EXU/CSRControl/_1681_ ( .A(\EXU/CSRControl/_0841_ ), .ZN(\EXU/CSRControl/_0842_ ) );
BUF_X4 \EXU/CSRControl/_1682_ ( .A(\EXU/CSRControl/_0842_ ), .Z(\EXU/CSRControl/_0843_ ) );
AOI211_X2 \EXU/CSRControl/_1683_ ( .A(\EXU/CSRControl/_0798_ ), .B(\EXU/CSRControl/_0802_ ), .C1(\EXU/CSRControl/_0839_ ), .C2(\EXU/CSRControl/_0843_ ), .ZN(\EXU/CSRControl/_0307_ ) );
NOR4_X1 \EXU/CSRControl/_1684_ ( .A1(\EXU/CSRControl/_0801_ ), .A2(fanout_net_18 ), .A3(fanout_net_17 ), .A4(\EXU/CSRControl/_0175_ ), .ZN(\EXU/CSRControl/_0844_ ) );
NAND3_X1 \EXU/CSRControl/_1685_ ( .A1(\EXU/CSRControl/_0813_ ), .A2(\EXU/CSRControl/_0175_ ), .A3(\EXU/CSRControl/_0816_ ), .ZN(\EXU/CSRControl/_0845_ ) );
BUF_X4 \EXU/CSRControl/_1686_ ( .A(\EXU/CSRControl/_0815_ ), .Z(\EXU/CSRControl/_0846_ ) );
NAND3_X1 \EXU/CSRControl/_1687_ ( .A1(\EXU/CSRControl/_0821_ ), .A2(\EXU/CSRControl/_0239_ ), .A3(\EXU/CSRControl/_0846_ ), .ZN(\EXU/CSRControl/_0847_ ) );
NAND4_X1 \EXU/CSRControl/_1688_ ( .A1(\EXU/CSRControl/_0827_ ), .A2(\EXU/CSRControl/_0829_ ), .A3(\EXU/CSRControl/_0207_ ), .A4(\EXU/CSRControl/_0830_ ), .ZN(\EXU/CSRControl/_0848_ ) );
AND3_X1 \EXU/CSRControl/_1689_ ( .A1(\EXU/CSRControl/_0845_ ), .A2(\EXU/CSRControl/_0847_ ), .A3(\EXU/CSRControl/_0848_ ), .ZN(\EXU/CSRControl/_0849_ ) );
NAND3_X1 \EXU/CSRControl/_1690_ ( .A1(\EXU/CSRControl/_0834_ ), .A2(\EXU/CSRControl/_0143_ ), .A3(\EXU/CSRControl/_0835_ ), .ZN(\EXU/CSRControl/_0850_ ) );
AOI21_X1 \EXU/CSRControl/_1691_ ( .A(\EXU/CSRControl/_0805_ ), .B1(\EXU/CSRControl/_0849_ ), .B2(\EXU/CSRControl/_0850_ ), .ZN(\EXU/CSRControl/_0851_ ) );
AOI21_X1 \EXU/CSRControl/_1692_ ( .A(\EXU/CSRControl/_0851_ ), .B1(\EXU/CSRControl/_0207_ ), .B2(\EXU/CSRControl/_0838_ ), .ZN(\EXU/CSRControl/_0852_ ) );
AOI211_X2 \EXU/CSRControl/_1693_ ( .A(\EXU/CSRControl/_0798_ ), .B(\EXU/CSRControl/_0844_ ), .C1(\EXU/CSRControl/_0852_ ), .C2(\EXU/CSRControl/_0843_ ), .ZN(\EXU/CSRControl/_0318_ ) );
NOR4_X1 \EXU/CSRControl/_1694_ ( .A1(\EXU/CSRControl/_0801_ ), .A2(fanout_net_18 ), .A3(fanout_net_17 ), .A4(\EXU/CSRControl/_0186_ ), .ZN(\EXU/CSRControl/_0853_ ) );
NAND3_X1 \EXU/CSRControl/_1695_ ( .A1(\EXU/CSRControl/_0813_ ), .A2(\EXU/CSRControl/_0186_ ), .A3(\EXU/CSRControl/_0816_ ), .ZN(\EXU/CSRControl/_0854_ ) );
NAND3_X1 \EXU/CSRControl/_1696_ ( .A1(\EXU/CSRControl/_0821_ ), .A2(\EXU/CSRControl/_0250_ ), .A3(\EXU/CSRControl/_0846_ ), .ZN(\EXU/CSRControl/_0855_ ) );
NAND4_X1 \EXU/CSRControl/_1697_ ( .A1(\EXU/CSRControl/_0827_ ), .A2(\EXU/CSRControl/_0829_ ), .A3(\EXU/CSRControl/_0218_ ), .A4(\EXU/CSRControl/_0830_ ), .ZN(\EXU/CSRControl/_0856_ ) );
AND3_X1 \EXU/CSRControl/_1698_ ( .A1(\EXU/CSRControl/_0854_ ), .A2(\EXU/CSRControl/_0855_ ), .A3(\EXU/CSRControl/_0856_ ), .ZN(\EXU/CSRControl/_0857_ ) );
NAND3_X1 \EXU/CSRControl/_1699_ ( .A1(\EXU/CSRControl/_0834_ ), .A2(\EXU/CSRControl/_0154_ ), .A3(\EXU/CSRControl/_0835_ ), .ZN(\EXU/CSRControl/_0858_ ) );
AOI21_X1 \EXU/CSRControl/_1700_ ( .A(\EXU/CSRControl/_0805_ ), .B1(\EXU/CSRControl/_0857_ ), .B2(\EXU/CSRControl/_0858_ ), .ZN(\EXU/CSRControl/_0859_ ) );
AOI21_X1 \EXU/CSRControl/_1701_ ( .A(\EXU/CSRControl/_0859_ ), .B1(\EXU/CSRControl/_0218_ ), .B2(\EXU/CSRControl/_0838_ ), .ZN(\EXU/CSRControl/_0860_ ) );
AOI211_X2 \EXU/CSRControl/_1702_ ( .A(\EXU/CSRControl/_0798_ ), .B(\EXU/CSRControl/_0853_ ), .C1(\EXU/CSRControl/_0860_ ), .C2(\EXU/CSRControl/_0843_ ), .ZN(\EXU/CSRControl/_0329_ ) );
NOR4_X1 \EXU/CSRControl/_1703_ ( .A1(\EXU/CSRControl/_0801_ ), .A2(fanout_net_18 ), .A3(fanout_net_17 ), .A4(\EXU/CSRControl/_0189_ ), .ZN(\EXU/CSRControl/_0861_ ) );
INV_X16 \EXU/CSRControl/_1704_ ( .A(\EXU/CSRControl/_0267_ ), .ZN(\EXU/CSRControl/_0862_ ) );
NAND4_X1 \EXU/CSRControl/_1705_ ( .A1(\EXU/CSRControl/_0828_ ), .A2(\EXU/CSRControl/_0862_ ), .A3(\EXU/CSRControl/_0266_ ), .A4(\EXU/CSRControl/_0808_ ), .ZN(\EXU/CSRControl/_0863_ ) );
NAND4_X1 \EXU/CSRControl/_1706_ ( .A1(\EXU/CSRControl/_0271_ ), .A2(\EXU/CSRControl/_0270_ ), .A3(\EXU/CSRControl/_0262_ ), .A4(\EXU/CSRControl/_0261_ ), .ZN(\EXU/CSRControl/_0864_ ) );
NOR2_X2 \EXU/CSRControl/_1707_ ( .A1(\EXU/CSRControl/_0863_ ), .A2(\EXU/CSRControl/_0864_ ), .ZN(\EXU/CSRControl/_0865_ ) );
INV_X1 \EXU/CSRControl/_1708_ ( .A(\EXU/CSRControl/_0865_ ), .ZN(\EXU/CSRControl/_0866_ ) );
CLKBUF_X2 \EXU/CSRControl/_1709_ ( .A(\EXU/CSRControl/_0866_ ), .Z(\EXU/CSRControl/_0867_ ) );
BUF_X8 \EXU/CSRControl/_1710_ ( .A(\EXU/CSRControl/_0812_ ), .Z(\EXU/CSRControl/_0868_ ) );
BUF_X2 \EXU/CSRControl/_1711_ ( .A(\EXU/CSRControl/_0815_ ), .Z(\EXU/CSRControl/_0869_ ) );
NAND3_X1 \EXU/CSRControl/_1712_ ( .A1(\EXU/CSRControl/_0868_ ), .A2(\EXU/CSRControl/_0189_ ), .A3(\EXU/CSRControl/_0869_ ), .ZN(\EXU/CSRControl/_0870_ ) );
BUF_X4 \EXU/CSRControl/_1713_ ( .A(\EXU/CSRControl/_0820_ ), .Z(\EXU/CSRControl/_0871_ ) );
BUF_X4 \EXU/CSRControl/_1714_ ( .A(\EXU/CSRControl/_0815_ ), .Z(\EXU/CSRControl/_0872_ ) );
NAND3_X1 \EXU/CSRControl/_1715_ ( .A1(\EXU/CSRControl/_0871_ ), .A2(\EXU/CSRControl/_0253_ ), .A3(\EXU/CSRControl/_0872_ ), .ZN(\EXU/CSRControl/_0873_ ) );
BUF_X4 \EXU/CSRControl/_1716_ ( .A(\EXU/CSRControl/_0826_ ), .Z(\EXU/CSRControl/_0874_ ) );
BUF_X4 \EXU/CSRControl/_1717_ ( .A(\EXU/CSRControl/_0828_ ), .Z(\EXU/CSRControl/_0875_ ) );
BUF_X4 \EXU/CSRControl/_1718_ ( .A(\EXU/CSRControl/_0815_ ), .Z(\EXU/CSRControl/_0876_ ) );
NAND4_X1 \EXU/CSRControl/_1719_ ( .A1(\EXU/CSRControl/_0874_ ), .A2(\EXU/CSRControl/_0875_ ), .A3(\EXU/CSRControl/_0221_ ), .A4(\EXU/CSRControl/_0876_ ), .ZN(\EXU/CSRControl/_0877_ ) );
AND4_X1 \EXU/CSRControl/_1720_ ( .A1(\EXU/CSRControl/_0867_ ), .A2(\EXU/CSRControl/_0870_ ), .A3(\EXU/CSRControl/_0873_ ), .A4(\EXU/CSRControl/_0877_ ), .ZN(\EXU/CSRControl/_0878_ ) );
NAND3_X1 \EXU/CSRControl/_1721_ ( .A1(\EXU/CSRControl/_0834_ ), .A2(\EXU/CSRControl/_0157_ ), .A3(\EXU/CSRControl/_0835_ ), .ZN(\EXU/CSRControl/_0879_ ) );
AOI21_X1 \EXU/CSRControl/_1722_ ( .A(\EXU/CSRControl/_0805_ ), .B1(\EXU/CSRControl/_0878_ ), .B2(\EXU/CSRControl/_0879_ ), .ZN(\EXU/CSRControl/_0880_ ) );
AOI21_X1 \EXU/CSRControl/_1723_ ( .A(\EXU/CSRControl/_0880_ ), .B1(\EXU/CSRControl/_0221_ ), .B2(\EXU/CSRControl/_0838_ ), .ZN(\EXU/CSRControl/_0881_ ) );
AOI211_X2 \EXU/CSRControl/_1724_ ( .A(\EXU/CSRControl/_0798_ ), .B(\EXU/CSRControl/_0861_ ), .C1(\EXU/CSRControl/_0881_ ), .C2(\EXU/CSRControl/_0843_ ), .ZN(\EXU/CSRControl/_0332_ ) );
NOR4_X1 \EXU/CSRControl/_1725_ ( .A1(\EXU/CSRControl/_0801_ ), .A2(fanout_net_18 ), .A3(fanout_net_17 ), .A4(\EXU/CSRControl/_0190_ ), .ZN(\EXU/CSRControl/_0882_ ) );
BUF_X4 \EXU/CSRControl/_1726_ ( .A(\EXU/CSRControl/_0804_ ), .Z(\EXU/CSRControl/_0883_ ) );
BUF_X4 \EXU/CSRControl/_1727_ ( .A(\EXU/CSRControl/_0883_ ), .Z(\EXU/CSRControl/_0884_ ) );
NAND3_X1 \EXU/CSRControl/_1728_ ( .A1(\EXU/CSRControl/_0868_ ), .A2(\EXU/CSRControl/_0190_ ), .A3(\EXU/CSRControl/_0869_ ), .ZN(\EXU/CSRControl/_0885_ ) );
NAND3_X1 \EXU/CSRControl/_1729_ ( .A1(\EXU/CSRControl/_0871_ ), .A2(\EXU/CSRControl/_0254_ ), .A3(\EXU/CSRControl/_0872_ ), .ZN(\EXU/CSRControl/_0886_ ) );
NAND4_X1 \EXU/CSRControl/_1730_ ( .A1(\EXU/CSRControl/_0874_ ), .A2(\EXU/CSRControl/_0875_ ), .A3(\EXU/CSRControl/_0222_ ), .A4(\EXU/CSRControl/_0876_ ), .ZN(\EXU/CSRControl/_0887_ ) );
AND4_X1 \EXU/CSRControl/_1731_ ( .A1(\EXU/CSRControl/_0867_ ), .A2(\EXU/CSRControl/_0885_ ), .A3(\EXU/CSRControl/_0886_ ), .A4(\EXU/CSRControl/_0887_ ), .ZN(\EXU/CSRControl/_0888_ ) );
NAND3_X1 \EXU/CSRControl/_1732_ ( .A1(\EXU/CSRControl/_0834_ ), .A2(\EXU/CSRControl/_0158_ ), .A3(\EXU/CSRControl/_0835_ ), .ZN(\EXU/CSRControl/_0889_ ) );
AOI21_X1 \EXU/CSRControl/_1733_ ( .A(\EXU/CSRControl/_0884_ ), .B1(\EXU/CSRControl/_0888_ ), .B2(\EXU/CSRControl/_0889_ ), .ZN(\EXU/CSRControl/_0890_ ) );
AOI21_X1 \EXU/CSRControl/_1734_ ( .A(\EXU/CSRControl/_0890_ ), .B1(\EXU/CSRControl/_0222_ ), .B2(\EXU/CSRControl/_0838_ ), .ZN(\EXU/CSRControl/_0891_ ) );
AOI211_X2 \EXU/CSRControl/_1735_ ( .A(\EXU/CSRControl/_0798_ ), .B(\EXU/CSRControl/_0882_ ), .C1(\EXU/CSRControl/_0891_ ), .C2(\EXU/CSRControl/_0843_ ), .ZN(\EXU/CSRControl/_0333_ ) );
NOR4_X1 \EXU/CSRControl/_1736_ ( .A1(\EXU/CSRControl/_0801_ ), .A2(fanout_net_18 ), .A3(fanout_net_17 ), .A4(\EXU/CSRControl/_0191_ ), .ZN(\EXU/CSRControl/_0892_ ) );
NAND3_X1 \EXU/CSRControl/_1737_ ( .A1(\EXU/CSRControl/_0868_ ), .A2(\EXU/CSRControl/_0191_ ), .A3(\EXU/CSRControl/_0869_ ), .ZN(\EXU/CSRControl/_0893_ ) );
NAND3_X1 \EXU/CSRControl/_1738_ ( .A1(\EXU/CSRControl/_0871_ ), .A2(\EXU/CSRControl/_0255_ ), .A3(\EXU/CSRControl/_0872_ ), .ZN(\EXU/CSRControl/_0894_ ) );
NAND4_X1 \EXU/CSRControl/_1739_ ( .A1(\EXU/CSRControl/_0874_ ), .A2(\EXU/CSRControl/_0875_ ), .A3(\EXU/CSRControl/_0223_ ), .A4(\EXU/CSRControl/_0876_ ), .ZN(\EXU/CSRControl/_0895_ ) );
AND4_X1 \EXU/CSRControl/_1740_ ( .A1(\EXU/CSRControl/_0867_ ), .A2(\EXU/CSRControl/_0893_ ), .A3(\EXU/CSRControl/_0894_ ), .A4(\EXU/CSRControl/_0895_ ), .ZN(\EXU/CSRControl/_0896_ ) );
NAND3_X1 \EXU/CSRControl/_1741_ ( .A1(\EXU/CSRControl/_0834_ ), .A2(\EXU/CSRControl/_0159_ ), .A3(\EXU/CSRControl/_0835_ ), .ZN(\EXU/CSRControl/_0897_ ) );
AOI21_X1 \EXU/CSRControl/_1742_ ( .A(\EXU/CSRControl/_0884_ ), .B1(\EXU/CSRControl/_0896_ ), .B2(\EXU/CSRControl/_0897_ ), .ZN(\EXU/CSRControl/_0898_ ) );
AOI21_X1 \EXU/CSRControl/_1743_ ( .A(\EXU/CSRControl/_0898_ ), .B1(\EXU/CSRControl/_0223_ ), .B2(\EXU/CSRControl/_0838_ ), .ZN(\EXU/CSRControl/_0899_ ) );
AOI211_X2 \EXU/CSRControl/_1744_ ( .A(\EXU/CSRControl/_0798_ ), .B(\EXU/CSRControl/_0892_ ), .C1(\EXU/CSRControl/_0899_ ), .C2(\EXU/CSRControl/_0843_ ), .ZN(\EXU/CSRControl/_0334_ ) );
NOR4_X1 \EXU/CSRControl/_1745_ ( .A1(\EXU/CSRControl/_0801_ ), .A2(fanout_net_18 ), .A3(fanout_net_17 ), .A4(\EXU/CSRControl/_0192_ ), .ZN(\EXU/CSRControl/_0900_ ) );
NAND3_X1 \EXU/CSRControl/_1746_ ( .A1(\EXU/CSRControl/_0868_ ), .A2(\EXU/CSRControl/_0192_ ), .A3(\EXU/CSRControl/_0822_ ), .ZN(\EXU/CSRControl/_0901_ ) );
NAND3_X1 \EXU/CSRControl/_1747_ ( .A1(\EXU/CSRControl/_0871_ ), .A2(\EXU/CSRControl/_0256_ ), .A3(\EXU/CSRControl/_0869_ ), .ZN(\EXU/CSRControl/_0902_ ) );
BUF_X4 \EXU/CSRControl/_1748_ ( .A(\EXU/CSRControl/_0826_ ), .Z(\EXU/CSRControl/_0903_ ) );
NAND4_X1 \EXU/CSRControl/_1749_ ( .A1(\EXU/CSRControl/_0903_ ), .A2(\EXU/CSRControl/_0875_ ), .A3(\EXU/CSRControl/_0224_ ), .A4(\EXU/CSRControl/_0872_ ), .ZN(\EXU/CSRControl/_0904_ ) );
NAND3_X1 \EXU/CSRControl/_1750_ ( .A1(\EXU/CSRControl/_0901_ ), .A2(\EXU/CSRControl/_0902_ ), .A3(\EXU/CSRControl/_0904_ ), .ZN(\EXU/CSRControl/_0905_ ) );
NOR2_X1 \EXU/CSRControl/_1751_ ( .A1(\EXU/CSRControl/_0905_ ), .A2(\EXU/CSRControl/_0865_ ), .ZN(\EXU/CSRControl/_0906_ ) );
NAND3_X1 \EXU/CSRControl/_1752_ ( .A1(\EXU/CSRControl/_0834_ ), .A2(\EXU/CSRControl/_0160_ ), .A3(\EXU/CSRControl/_0835_ ), .ZN(\EXU/CSRControl/_0907_ ) );
AOI21_X1 \EXU/CSRControl/_1753_ ( .A(\EXU/CSRControl/_0884_ ), .B1(\EXU/CSRControl/_0906_ ), .B2(\EXU/CSRControl/_0907_ ), .ZN(\EXU/CSRControl/_0908_ ) );
AOI21_X1 \EXU/CSRControl/_1754_ ( .A(\EXU/CSRControl/_0908_ ), .B1(\EXU/CSRControl/_0224_ ), .B2(\EXU/CSRControl/_0838_ ), .ZN(\EXU/CSRControl/_0909_ ) );
AOI211_X2 \EXU/CSRControl/_1755_ ( .A(\EXU/CSRControl/_0798_ ), .B(\EXU/CSRControl/_0900_ ), .C1(\EXU/CSRControl/_0909_ ), .C2(\EXU/CSRControl/_0843_ ), .ZN(\EXU/CSRControl/_0335_ ) );
NOR4_X1 \EXU/CSRControl/_1756_ ( .A1(\EXU/CSRControl/_0801_ ), .A2(fanout_net_18 ), .A3(fanout_net_17 ), .A4(\EXU/CSRControl/_0193_ ), .ZN(\EXU/CSRControl/_0910_ ) );
NAND3_X1 \EXU/CSRControl/_1757_ ( .A1(\EXU/CSRControl/_0813_ ), .A2(\EXU/CSRControl/_0193_ ), .A3(\EXU/CSRControl/_0816_ ), .ZN(\EXU/CSRControl/_0911_ ) );
NAND3_X1 \EXU/CSRControl/_1758_ ( .A1(\EXU/CSRControl/_0821_ ), .A2(\EXU/CSRControl/_0257_ ), .A3(\EXU/CSRControl/_0846_ ), .ZN(\EXU/CSRControl/_0912_ ) );
NAND4_X1 \EXU/CSRControl/_1759_ ( .A1(\EXU/CSRControl/_0827_ ), .A2(\EXU/CSRControl/_0829_ ), .A3(\EXU/CSRControl/_0225_ ), .A4(\EXU/CSRControl/_0830_ ), .ZN(\EXU/CSRControl/_0913_ ) );
AND3_X1 \EXU/CSRControl/_1760_ ( .A1(\EXU/CSRControl/_0911_ ), .A2(\EXU/CSRControl/_0912_ ), .A3(\EXU/CSRControl/_0913_ ), .ZN(\EXU/CSRControl/_0914_ ) );
NAND3_X1 \EXU/CSRControl/_1761_ ( .A1(\EXU/CSRControl/_0834_ ), .A2(\EXU/CSRControl/_0161_ ), .A3(\EXU/CSRControl/_0835_ ), .ZN(\EXU/CSRControl/_0915_ ) );
AOI21_X1 \EXU/CSRControl/_1762_ ( .A(\EXU/CSRControl/_0884_ ), .B1(\EXU/CSRControl/_0914_ ), .B2(\EXU/CSRControl/_0915_ ), .ZN(\EXU/CSRControl/_0916_ ) );
AOI21_X1 \EXU/CSRControl/_1763_ ( .A(\EXU/CSRControl/_0916_ ), .B1(\EXU/CSRControl/_0225_ ), .B2(\EXU/CSRControl/_0838_ ), .ZN(\EXU/CSRControl/_0917_ ) );
AOI211_X2 \EXU/CSRControl/_1764_ ( .A(\EXU/CSRControl/_0798_ ), .B(\EXU/CSRControl/_0910_ ), .C1(\EXU/CSRControl/_0917_ ), .C2(\EXU/CSRControl/_0843_ ), .ZN(\EXU/CSRControl/_0336_ ) );
NOR4_X1 \EXU/CSRControl/_1765_ ( .A1(\EXU/CSRControl/_0801_ ), .A2(fanout_net_18 ), .A3(fanout_net_17 ), .A4(\EXU/CSRControl/_0194_ ), .ZN(\EXU/CSRControl/_0918_ ) );
NAND3_X1 \EXU/CSRControl/_1766_ ( .A1(\EXU/CSRControl/_0868_ ), .A2(\EXU/CSRControl/_0194_ ), .A3(\EXU/CSRControl/_0869_ ), .ZN(\EXU/CSRControl/_0919_ ) );
NAND3_X1 \EXU/CSRControl/_1767_ ( .A1(\EXU/CSRControl/_0871_ ), .A2(\EXU/CSRControl/_0258_ ), .A3(\EXU/CSRControl/_0872_ ), .ZN(\EXU/CSRControl/_0920_ ) );
NAND4_X1 \EXU/CSRControl/_1768_ ( .A1(\EXU/CSRControl/_0874_ ), .A2(\EXU/CSRControl/_0875_ ), .A3(\EXU/CSRControl/_0226_ ), .A4(\EXU/CSRControl/_0876_ ), .ZN(\EXU/CSRControl/_0921_ ) );
AND4_X1 \EXU/CSRControl/_1769_ ( .A1(\EXU/CSRControl/_0867_ ), .A2(\EXU/CSRControl/_0919_ ), .A3(\EXU/CSRControl/_0920_ ), .A4(\EXU/CSRControl/_0921_ ), .ZN(\EXU/CSRControl/_0922_ ) );
NAND3_X1 \EXU/CSRControl/_1770_ ( .A1(\EXU/CSRControl/_0834_ ), .A2(\EXU/CSRControl/_0162_ ), .A3(\EXU/CSRControl/_0835_ ), .ZN(\EXU/CSRControl/_0923_ ) );
AOI21_X1 \EXU/CSRControl/_1771_ ( .A(\EXU/CSRControl/_0884_ ), .B1(\EXU/CSRControl/_0922_ ), .B2(\EXU/CSRControl/_0923_ ), .ZN(\EXU/CSRControl/_0924_ ) );
AOI21_X1 \EXU/CSRControl/_1772_ ( .A(\EXU/CSRControl/_0924_ ), .B1(\EXU/CSRControl/_0226_ ), .B2(\EXU/CSRControl/_0838_ ), .ZN(\EXU/CSRControl/_0925_ ) );
AOI211_X2 \EXU/CSRControl/_1773_ ( .A(\EXU/CSRControl/_0798_ ), .B(\EXU/CSRControl/_0918_ ), .C1(\EXU/CSRControl/_0925_ ), .C2(\EXU/CSRControl/_0843_ ), .ZN(\EXU/CSRControl/_0337_ ) );
BUF_X4 \EXU/CSRControl/_1774_ ( .A(\EXU/CSRControl/_0800_ ), .Z(\EXU/CSRControl/_0926_ ) );
NOR4_X1 \EXU/CSRControl/_1775_ ( .A1(\EXU/CSRControl/_0926_ ), .A2(fanout_net_18 ), .A3(fanout_net_17 ), .A4(\EXU/CSRControl/_0195_ ), .ZN(\EXU/CSRControl/_0927_ ) );
NAND3_X1 \EXU/CSRControl/_1776_ ( .A1(\EXU/CSRControl/_0813_ ), .A2(\EXU/CSRControl/_0195_ ), .A3(\EXU/CSRControl/_0816_ ), .ZN(\EXU/CSRControl/_0928_ ) );
NAND3_X1 \EXU/CSRControl/_1777_ ( .A1(\EXU/CSRControl/_0821_ ), .A2(\EXU/CSRControl/_0259_ ), .A3(\EXU/CSRControl/_0846_ ), .ZN(\EXU/CSRControl/_0929_ ) );
NAND4_X1 \EXU/CSRControl/_1778_ ( .A1(\EXU/CSRControl/_0903_ ), .A2(\EXU/CSRControl/_0829_ ), .A3(\EXU/CSRControl/_0227_ ), .A4(\EXU/CSRControl/_0830_ ), .ZN(\EXU/CSRControl/_0930_ ) );
AND3_X1 \EXU/CSRControl/_1779_ ( .A1(\EXU/CSRControl/_0928_ ), .A2(\EXU/CSRControl/_0929_ ), .A3(\EXU/CSRControl/_0930_ ), .ZN(\EXU/CSRControl/_0931_ ) );
NAND3_X1 \EXU/CSRControl/_1780_ ( .A1(\EXU/CSRControl/_0834_ ), .A2(\EXU/CSRControl/_0163_ ), .A3(\EXU/CSRControl/_0835_ ), .ZN(\EXU/CSRControl/_0932_ ) );
AOI21_X1 \EXU/CSRControl/_1781_ ( .A(\EXU/CSRControl/_0884_ ), .B1(\EXU/CSRControl/_0931_ ), .B2(\EXU/CSRControl/_0932_ ), .ZN(\EXU/CSRControl/_0933_ ) );
AOI21_X1 \EXU/CSRControl/_1782_ ( .A(\EXU/CSRControl/_0933_ ), .B1(\EXU/CSRControl/_0227_ ), .B2(\EXU/CSRControl/_0838_ ), .ZN(\EXU/CSRControl/_0934_ ) );
BUF_X4 \EXU/CSRControl/_1783_ ( .A(\EXU/CSRControl/_0842_ ), .Z(\EXU/CSRControl/_0935_ ) );
AOI211_X2 \EXU/CSRControl/_1784_ ( .A(\EXU/CSRControl/_0798_ ), .B(\EXU/CSRControl/_0927_ ), .C1(\EXU/CSRControl/_0934_ ), .C2(\EXU/CSRControl/_0935_ ), .ZN(\EXU/CSRControl/_0338_ ) );
BUF_X4 \EXU/CSRControl/_1785_ ( .A(\EXU/CSRControl/_0797_ ), .Z(\EXU/CSRControl/_0936_ ) );
NOR4_X1 \EXU/CSRControl/_1786_ ( .A1(\EXU/CSRControl/_0926_ ), .A2(fanout_net_18 ), .A3(fanout_net_17 ), .A4(\EXU/CSRControl/_0165_ ), .ZN(\EXU/CSRControl/_0937_ ) );
NAND3_X1 \EXU/CSRControl/_1787_ ( .A1(\EXU/CSRControl/_0813_ ), .A2(\EXU/CSRControl/_0165_ ), .A3(\EXU/CSRControl/_0822_ ), .ZN(\EXU/CSRControl/_0938_ ) );
NAND3_X1 \EXU/CSRControl/_1788_ ( .A1(\EXU/CSRControl/_0821_ ), .A2(\EXU/CSRControl/_0229_ ), .A3(\EXU/CSRControl/_0846_ ), .ZN(\EXU/CSRControl/_0939_ ) );
NAND4_X1 \EXU/CSRControl/_1789_ ( .A1(\EXU/CSRControl/_0903_ ), .A2(\EXU/CSRControl/_0829_ ), .A3(\EXU/CSRControl/_0197_ ), .A4(\EXU/CSRControl/_0830_ ), .ZN(\EXU/CSRControl/_0940_ ) );
AND3_X1 \EXU/CSRControl/_1790_ ( .A1(\EXU/CSRControl/_0938_ ), .A2(\EXU/CSRControl/_0939_ ), .A3(\EXU/CSRControl/_0940_ ), .ZN(\EXU/CSRControl/_0941_ ) );
BUF_X4 \EXU/CSRControl/_1791_ ( .A(\EXU/CSRControl/_0833_ ), .Z(\EXU/CSRControl/_0942_ ) );
BUF_X4 \EXU/CSRControl/_1792_ ( .A(\EXU/CSRControl/_0816_ ), .Z(\EXU/CSRControl/_0943_ ) );
NAND3_X1 \EXU/CSRControl/_1793_ ( .A1(\EXU/CSRControl/_0942_ ), .A2(\EXU/CSRControl/_0133_ ), .A3(\EXU/CSRControl/_0943_ ), .ZN(\EXU/CSRControl/_0944_ ) );
AOI21_X1 \EXU/CSRControl/_1794_ ( .A(\EXU/CSRControl/_0884_ ), .B1(\EXU/CSRControl/_0941_ ), .B2(\EXU/CSRControl/_0944_ ), .ZN(\EXU/CSRControl/_0945_ ) );
BUF_X4 \EXU/CSRControl/_1795_ ( .A(\EXU/CSRControl/_0805_ ), .Z(\EXU/CSRControl/_0946_ ) );
AOI21_X1 \EXU/CSRControl/_1796_ ( .A(\EXU/CSRControl/_0945_ ), .B1(\EXU/CSRControl/_0197_ ), .B2(\EXU/CSRControl/_0946_ ), .ZN(\EXU/CSRControl/_0947_ ) );
AOI211_X2 \EXU/CSRControl/_1797_ ( .A(\EXU/CSRControl/_0936_ ), .B(\EXU/CSRControl/_0937_ ), .C1(\EXU/CSRControl/_0947_ ), .C2(\EXU/CSRControl/_0935_ ), .ZN(\EXU/CSRControl/_0308_ ) );
NOR4_X1 \EXU/CSRControl/_1798_ ( .A1(\EXU/CSRControl/_0926_ ), .A2(fanout_net_18 ), .A3(fanout_net_17 ), .A4(\EXU/CSRControl/_0166_ ), .ZN(\EXU/CSRControl/_0948_ ) );
NAND3_X1 \EXU/CSRControl/_1799_ ( .A1(\EXU/CSRControl/_0868_ ), .A2(\EXU/CSRControl/_0166_ ), .A3(\EXU/CSRControl/_0869_ ), .ZN(\EXU/CSRControl/_0949_ ) );
NAND3_X1 \EXU/CSRControl/_1800_ ( .A1(\EXU/CSRControl/_0871_ ), .A2(\EXU/CSRControl/_0230_ ), .A3(\EXU/CSRControl/_0872_ ), .ZN(\EXU/CSRControl/_0950_ ) );
NAND4_X1 \EXU/CSRControl/_1801_ ( .A1(\EXU/CSRControl/_0874_ ), .A2(\EXU/CSRControl/_0875_ ), .A3(\EXU/CSRControl/_0198_ ), .A4(\EXU/CSRControl/_0876_ ), .ZN(\EXU/CSRControl/_0951_ ) );
AND4_X1 \EXU/CSRControl/_1802_ ( .A1(\EXU/CSRControl/_0867_ ), .A2(\EXU/CSRControl/_0949_ ), .A3(\EXU/CSRControl/_0950_ ), .A4(\EXU/CSRControl/_0951_ ), .ZN(\EXU/CSRControl/_0952_ ) );
NAND3_X1 \EXU/CSRControl/_1803_ ( .A1(\EXU/CSRControl/_0942_ ), .A2(\EXU/CSRControl/_0134_ ), .A3(\EXU/CSRControl/_0943_ ), .ZN(\EXU/CSRControl/_0953_ ) );
AOI21_X1 \EXU/CSRControl/_1804_ ( .A(\EXU/CSRControl/_0884_ ), .B1(\EXU/CSRControl/_0952_ ), .B2(\EXU/CSRControl/_0953_ ), .ZN(\EXU/CSRControl/_0954_ ) );
AOI21_X1 \EXU/CSRControl/_1805_ ( .A(\EXU/CSRControl/_0954_ ), .B1(\EXU/CSRControl/_0198_ ), .B2(\EXU/CSRControl/_0946_ ), .ZN(\EXU/CSRControl/_0955_ ) );
AOI211_X2 \EXU/CSRControl/_1806_ ( .A(\EXU/CSRControl/_0936_ ), .B(\EXU/CSRControl/_0948_ ), .C1(\EXU/CSRControl/_0955_ ), .C2(\EXU/CSRControl/_0935_ ), .ZN(\EXU/CSRControl/_0309_ ) );
NOR4_X1 \EXU/CSRControl/_1807_ ( .A1(\EXU/CSRControl/_0926_ ), .A2(fanout_net_18 ), .A3(fanout_net_17 ), .A4(\EXU/CSRControl/_0167_ ), .ZN(\EXU/CSRControl/_0956_ ) );
BUF_X4 \EXU/CSRControl/_1808_ ( .A(\EXU/CSRControl/_0812_ ), .Z(\EXU/CSRControl/_0957_ ) );
BUF_X4 \EXU/CSRControl/_1809_ ( .A(\EXU/CSRControl/_0815_ ), .Z(\EXU/CSRControl/_0958_ ) );
NAND3_X1 \EXU/CSRControl/_1810_ ( .A1(\EXU/CSRControl/_0957_ ), .A2(\EXU/CSRControl/_0167_ ), .A3(\EXU/CSRControl/_0958_ ), .ZN(\EXU/CSRControl/_0959_ ) );
BUF_X4 \EXU/CSRControl/_1811_ ( .A(\EXU/CSRControl/_0815_ ), .Z(\EXU/CSRControl/_0960_ ) );
NAND3_X1 \EXU/CSRControl/_1812_ ( .A1(\EXU/CSRControl/_0871_ ), .A2(\EXU/CSRControl/_0231_ ), .A3(\EXU/CSRControl/_0960_ ), .ZN(\EXU/CSRControl/_0961_ ) );
NAND4_X1 \EXU/CSRControl/_1813_ ( .A1(\EXU/CSRControl/_0874_ ), .A2(\EXU/CSRControl/_0875_ ), .A3(\EXU/CSRControl/_0199_ ), .A4(\EXU/CSRControl/_0876_ ), .ZN(\EXU/CSRControl/_0962_ ) );
AND4_X1 \EXU/CSRControl/_1814_ ( .A1(\EXU/CSRControl/_0867_ ), .A2(\EXU/CSRControl/_0959_ ), .A3(\EXU/CSRControl/_0961_ ), .A4(\EXU/CSRControl/_0962_ ), .ZN(\EXU/CSRControl/_0963_ ) );
NAND3_X1 \EXU/CSRControl/_1815_ ( .A1(\EXU/CSRControl/_0942_ ), .A2(\EXU/CSRControl/_0135_ ), .A3(\EXU/CSRControl/_0943_ ), .ZN(\EXU/CSRControl/_0964_ ) );
AOI21_X1 \EXU/CSRControl/_1816_ ( .A(\EXU/CSRControl/_0884_ ), .B1(\EXU/CSRControl/_0963_ ), .B2(\EXU/CSRControl/_0964_ ), .ZN(\EXU/CSRControl/_0965_ ) );
AOI21_X1 \EXU/CSRControl/_1817_ ( .A(\EXU/CSRControl/_0965_ ), .B1(\EXU/CSRControl/_0199_ ), .B2(\EXU/CSRControl/_0946_ ), .ZN(\EXU/CSRControl/_0966_ ) );
AOI211_X2 \EXU/CSRControl/_1818_ ( .A(\EXU/CSRControl/_0936_ ), .B(\EXU/CSRControl/_0956_ ), .C1(\EXU/CSRControl/_0966_ ), .C2(\EXU/CSRControl/_0935_ ), .ZN(\EXU/CSRControl/_0310_ ) );
NOR4_X1 \EXU/CSRControl/_1819_ ( .A1(\EXU/CSRControl/_0926_ ), .A2(fanout_net_18 ), .A3(fanout_net_17 ), .A4(\EXU/CSRControl/_0168_ ), .ZN(\EXU/CSRControl/_0967_ ) );
NAND3_X1 \EXU/CSRControl/_1820_ ( .A1(\EXU/CSRControl/_0957_ ), .A2(\EXU/CSRControl/_0168_ ), .A3(\EXU/CSRControl/_0958_ ), .ZN(\EXU/CSRControl/_0968_ ) );
BUF_X4 \EXU/CSRControl/_1821_ ( .A(\EXU/CSRControl/_0820_ ), .Z(\EXU/CSRControl/_0969_ ) );
NAND3_X1 \EXU/CSRControl/_1822_ ( .A1(\EXU/CSRControl/_0969_ ), .A2(\EXU/CSRControl/_0232_ ), .A3(\EXU/CSRControl/_0960_ ), .ZN(\EXU/CSRControl/_0970_ ) );
BUF_X4 \EXU/CSRControl/_1823_ ( .A(\EXU/CSRControl/_0828_ ), .Z(\EXU/CSRControl/_0971_ ) );
NAND4_X1 \EXU/CSRControl/_1824_ ( .A1(\EXU/CSRControl/_0874_ ), .A2(\EXU/CSRControl/_0971_ ), .A3(\EXU/CSRControl/_0200_ ), .A4(\EXU/CSRControl/_0876_ ), .ZN(\EXU/CSRControl/_0972_ ) );
AND4_X1 \EXU/CSRControl/_1825_ ( .A1(\EXU/CSRControl/_0867_ ), .A2(\EXU/CSRControl/_0968_ ), .A3(\EXU/CSRControl/_0970_ ), .A4(\EXU/CSRControl/_0972_ ), .ZN(\EXU/CSRControl/_0973_ ) );
NAND3_X1 \EXU/CSRControl/_1826_ ( .A1(\EXU/CSRControl/_0942_ ), .A2(\EXU/CSRControl/_0136_ ), .A3(\EXU/CSRControl/_0943_ ), .ZN(\EXU/CSRControl/_0974_ ) );
AOI21_X1 \EXU/CSRControl/_1827_ ( .A(\EXU/CSRControl/_0884_ ), .B1(\EXU/CSRControl/_0973_ ), .B2(\EXU/CSRControl/_0974_ ), .ZN(\EXU/CSRControl/_0975_ ) );
AOI21_X1 \EXU/CSRControl/_1828_ ( .A(\EXU/CSRControl/_0975_ ), .B1(\EXU/CSRControl/_0200_ ), .B2(\EXU/CSRControl/_0946_ ), .ZN(\EXU/CSRControl/_0976_ ) );
AOI211_X2 \EXU/CSRControl/_1829_ ( .A(\EXU/CSRControl/_0936_ ), .B(\EXU/CSRControl/_0967_ ), .C1(\EXU/CSRControl/_0976_ ), .C2(\EXU/CSRControl/_0935_ ), .ZN(\EXU/CSRControl/_0311_ ) );
NOR4_X1 \EXU/CSRControl/_1830_ ( .A1(\EXU/CSRControl/_0926_ ), .A2(fanout_net_18 ), .A3(fanout_net_17 ), .A4(\EXU/CSRControl/_0169_ ), .ZN(\EXU/CSRControl/_0977_ ) );
BUF_X4 \EXU/CSRControl/_1831_ ( .A(\EXU/CSRControl/_0804_ ), .Z(\EXU/CSRControl/_0978_ ) );
NAND3_X1 \EXU/CSRControl/_1832_ ( .A1(\EXU/CSRControl/_0957_ ), .A2(\EXU/CSRControl/_0169_ ), .A3(\EXU/CSRControl/_0958_ ), .ZN(\EXU/CSRControl/_0979_ ) );
NAND3_X1 \EXU/CSRControl/_1833_ ( .A1(\EXU/CSRControl/_0969_ ), .A2(\EXU/CSRControl/_0233_ ), .A3(\EXU/CSRControl/_0960_ ), .ZN(\EXU/CSRControl/_0980_ ) );
BUF_X4 \EXU/CSRControl/_1834_ ( .A(\EXU/CSRControl/_0826_ ), .Z(\EXU/CSRControl/_0981_ ) );
BUF_X4 \EXU/CSRControl/_1835_ ( .A(\EXU/CSRControl/_0814_ ), .Z(\EXU/CSRControl/_0982_ ) );
NAND4_X1 \EXU/CSRControl/_1836_ ( .A1(\EXU/CSRControl/_0981_ ), .A2(\EXU/CSRControl/_0971_ ), .A3(\EXU/CSRControl/_0201_ ), .A4(\EXU/CSRControl/_0982_ ), .ZN(\EXU/CSRControl/_0983_ ) );
AND4_X1 \EXU/CSRControl/_1837_ ( .A1(\EXU/CSRControl/_0867_ ), .A2(\EXU/CSRControl/_0979_ ), .A3(\EXU/CSRControl/_0980_ ), .A4(\EXU/CSRControl/_0983_ ), .ZN(\EXU/CSRControl/_0984_ ) );
NAND3_X1 \EXU/CSRControl/_1838_ ( .A1(\EXU/CSRControl/_0942_ ), .A2(\EXU/CSRControl/_0137_ ), .A3(\EXU/CSRControl/_0943_ ), .ZN(\EXU/CSRControl/_0985_ ) );
AOI21_X1 \EXU/CSRControl/_1839_ ( .A(\EXU/CSRControl/_0978_ ), .B1(\EXU/CSRControl/_0984_ ), .B2(\EXU/CSRControl/_0985_ ), .ZN(\EXU/CSRControl/_0986_ ) );
AOI21_X1 \EXU/CSRControl/_1840_ ( .A(\EXU/CSRControl/_0986_ ), .B1(\EXU/CSRControl/_0201_ ), .B2(\EXU/CSRControl/_0946_ ), .ZN(\EXU/CSRControl/_0987_ ) );
AOI211_X2 \EXU/CSRControl/_1841_ ( .A(\EXU/CSRControl/_0936_ ), .B(\EXU/CSRControl/_0977_ ), .C1(\EXU/CSRControl/_0987_ ), .C2(\EXU/CSRControl/_0935_ ), .ZN(\EXU/CSRControl/_0312_ ) );
NOR4_X1 \EXU/CSRControl/_1842_ ( .A1(\EXU/CSRControl/_0926_ ), .A2(fanout_net_18 ), .A3(fanout_net_17 ), .A4(\EXU/CSRControl/_0170_ ), .ZN(\EXU/CSRControl/_0988_ ) );
NAND3_X1 \EXU/CSRControl/_1843_ ( .A1(\EXU/CSRControl/_0813_ ), .A2(\EXU/CSRControl/_0170_ ), .A3(\EXU/CSRControl/_0822_ ), .ZN(\EXU/CSRControl/_0989_ ) );
NAND3_X1 \EXU/CSRControl/_1844_ ( .A1(\EXU/CSRControl/_0821_ ), .A2(\EXU/CSRControl/_0234_ ), .A3(\EXU/CSRControl/_0846_ ), .ZN(\EXU/CSRControl/_0990_ ) );
NAND4_X1 \EXU/CSRControl/_1845_ ( .A1(\EXU/CSRControl/_0903_ ), .A2(\EXU/CSRControl/_0829_ ), .A3(\EXU/CSRControl/_0202_ ), .A4(\EXU/CSRControl/_0830_ ), .ZN(\EXU/CSRControl/_0991_ ) );
AND3_X1 \EXU/CSRControl/_1846_ ( .A1(\EXU/CSRControl/_0989_ ), .A2(\EXU/CSRControl/_0990_ ), .A3(\EXU/CSRControl/_0991_ ), .ZN(\EXU/CSRControl/_0992_ ) );
NAND3_X1 \EXU/CSRControl/_1847_ ( .A1(\EXU/CSRControl/_0942_ ), .A2(\EXU/CSRControl/_0138_ ), .A3(\EXU/CSRControl/_0943_ ), .ZN(\EXU/CSRControl/_0993_ ) );
AOI21_X1 \EXU/CSRControl/_1848_ ( .A(\EXU/CSRControl/_0978_ ), .B1(\EXU/CSRControl/_0992_ ), .B2(\EXU/CSRControl/_0993_ ), .ZN(\EXU/CSRControl/_0994_ ) );
AOI21_X1 \EXU/CSRControl/_1849_ ( .A(\EXU/CSRControl/_0994_ ), .B1(\EXU/CSRControl/_0202_ ), .B2(\EXU/CSRControl/_0946_ ), .ZN(\EXU/CSRControl/_0995_ ) );
AOI211_X2 \EXU/CSRControl/_1850_ ( .A(\EXU/CSRControl/_0936_ ), .B(\EXU/CSRControl/_0988_ ), .C1(\EXU/CSRControl/_0995_ ), .C2(\EXU/CSRControl/_0935_ ), .ZN(\EXU/CSRControl/_0313_ ) );
NOR4_X1 \EXU/CSRControl/_1851_ ( .A1(\EXU/CSRControl/_0926_ ), .A2(fanout_net_18 ), .A3(fanout_net_17 ), .A4(\EXU/CSRControl/_0171_ ), .ZN(\EXU/CSRControl/_0996_ ) );
NAND3_X1 \EXU/CSRControl/_1852_ ( .A1(\EXU/CSRControl/_0957_ ), .A2(\EXU/CSRControl/_0171_ ), .A3(\EXU/CSRControl/_0958_ ), .ZN(\EXU/CSRControl/_0997_ ) );
NAND3_X1 \EXU/CSRControl/_1853_ ( .A1(\EXU/CSRControl/_0969_ ), .A2(\EXU/CSRControl/_0235_ ), .A3(\EXU/CSRControl/_0960_ ), .ZN(\EXU/CSRControl/_0998_ ) );
NAND4_X1 \EXU/CSRControl/_1854_ ( .A1(\EXU/CSRControl/_0981_ ), .A2(\EXU/CSRControl/_0971_ ), .A3(\EXU/CSRControl/_0203_ ), .A4(\EXU/CSRControl/_0982_ ), .ZN(\EXU/CSRControl/_0999_ ) );
AND4_X1 \EXU/CSRControl/_1855_ ( .A1(\EXU/CSRControl/_0867_ ), .A2(\EXU/CSRControl/_0997_ ), .A3(\EXU/CSRControl/_0998_ ), .A4(\EXU/CSRControl/_0999_ ), .ZN(\EXU/CSRControl/_1000_ ) );
NAND3_X1 \EXU/CSRControl/_1856_ ( .A1(\EXU/CSRControl/_0942_ ), .A2(\EXU/CSRControl/_0139_ ), .A3(\EXU/CSRControl/_0943_ ), .ZN(\EXU/CSRControl/_1001_ ) );
AOI21_X1 \EXU/CSRControl/_1857_ ( .A(\EXU/CSRControl/_0978_ ), .B1(\EXU/CSRControl/_1000_ ), .B2(\EXU/CSRControl/_1001_ ), .ZN(\EXU/CSRControl/_1002_ ) );
AOI21_X1 \EXU/CSRControl/_1858_ ( .A(\EXU/CSRControl/_1002_ ), .B1(\EXU/CSRControl/_0203_ ), .B2(\EXU/CSRControl/_0946_ ), .ZN(\EXU/CSRControl/_1003_ ) );
AOI211_X2 \EXU/CSRControl/_1859_ ( .A(\EXU/CSRControl/_0936_ ), .B(\EXU/CSRControl/_0996_ ), .C1(\EXU/CSRControl/_1003_ ), .C2(\EXU/CSRControl/_0935_ ), .ZN(\EXU/CSRControl/_0314_ ) );
NOR4_X1 \EXU/CSRControl/_1860_ ( .A1(\EXU/CSRControl/_0926_ ), .A2(fanout_net_18 ), .A3(fanout_net_17 ), .A4(\EXU/CSRControl/_0172_ ), .ZN(\EXU/CSRControl/_1004_ ) );
NAND3_X1 \EXU/CSRControl/_1861_ ( .A1(\EXU/CSRControl/_0957_ ), .A2(\EXU/CSRControl/_0172_ ), .A3(\EXU/CSRControl/_0958_ ), .ZN(\EXU/CSRControl/_1005_ ) );
NAND3_X1 \EXU/CSRControl/_1862_ ( .A1(\EXU/CSRControl/_0969_ ), .A2(\EXU/CSRControl/_0236_ ), .A3(\EXU/CSRControl/_0960_ ), .ZN(\EXU/CSRControl/_1006_ ) );
NAND4_X1 \EXU/CSRControl/_1863_ ( .A1(\EXU/CSRControl/_0981_ ), .A2(\EXU/CSRControl/_0971_ ), .A3(\EXU/CSRControl/_0204_ ), .A4(\EXU/CSRControl/_0982_ ), .ZN(\EXU/CSRControl/_1007_ ) );
AND4_X1 \EXU/CSRControl/_1864_ ( .A1(\EXU/CSRControl/_0867_ ), .A2(\EXU/CSRControl/_1005_ ), .A3(\EXU/CSRControl/_1006_ ), .A4(\EXU/CSRControl/_1007_ ), .ZN(\EXU/CSRControl/_1008_ ) );
NAND3_X1 \EXU/CSRControl/_1865_ ( .A1(\EXU/CSRControl/_0942_ ), .A2(\EXU/CSRControl/_0140_ ), .A3(\EXU/CSRControl/_0943_ ), .ZN(\EXU/CSRControl/_1009_ ) );
AOI21_X1 \EXU/CSRControl/_1866_ ( .A(\EXU/CSRControl/_0978_ ), .B1(\EXU/CSRControl/_1008_ ), .B2(\EXU/CSRControl/_1009_ ), .ZN(\EXU/CSRControl/_1010_ ) );
AOI21_X1 \EXU/CSRControl/_1867_ ( .A(\EXU/CSRControl/_1010_ ), .B1(\EXU/CSRControl/_0204_ ), .B2(\EXU/CSRControl/_0946_ ), .ZN(\EXU/CSRControl/_1011_ ) );
AOI211_X2 \EXU/CSRControl/_1868_ ( .A(\EXU/CSRControl/_0936_ ), .B(\EXU/CSRControl/_1004_ ), .C1(\EXU/CSRControl/_1011_ ), .C2(\EXU/CSRControl/_0935_ ), .ZN(\EXU/CSRControl/_0315_ ) );
NOR4_X1 \EXU/CSRControl/_1869_ ( .A1(\EXU/CSRControl/_0926_ ), .A2(fanout_net_18 ), .A3(fanout_net_17 ), .A4(\EXU/CSRControl/_0173_ ), .ZN(\EXU/CSRControl/_1012_ ) );
AND3_X1 \EXU/CSRControl/_1870_ ( .A1(\EXU/CSRControl/_0868_ ), .A2(\EXU/CSRControl/_0173_ ), .A3(\EXU/CSRControl/_0822_ ), .ZN(\EXU/CSRControl/_1013_ ) );
NAND4_X1 \EXU/CSRControl/_1871_ ( .A1(\EXU/CSRControl/_0827_ ), .A2(\EXU/CSRControl/_0829_ ), .A3(\EXU/CSRControl/_0205_ ), .A4(\EXU/CSRControl/_0869_ ), .ZN(\EXU/CSRControl/_1014_ ) );
NAND3_X1 \EXU/CSRControl/_1872_ ( .A1(\EXU/CSRControl/_0871_ ), .A2(\EXU/CSRControl/_0237_ ), .A3(\EXU/CSRControl/_0869_ ), .ZN(\EXU/CSRControl/_1015_ ) );
NAND2_X1 \EXU/CSRControl/_1873_ ( .A1(\EXU/CSRControl/_1014_ ), .A2(\EXU/CSRControl/_1015_ ), .ZN(\EXU/CSRControl/_1016_ ) );
NOR2_X1 \EXU/CSRControl/_1874_ ( .A1(\EXU/CSRControl/_1013_ ), .A2(\EXU/CSRControl/_1016_ ), .ZN(\EXU/CSRControl/_1017_ ) );
NAND3_X1 \EXU/CSRControl/_1875_ ( .A1(\EXU/CSRControl/_0942_ ), .A2(\EXU/CSRControl/_0141_ ), .A3(\EXU/CSRControl/_0943_ ), .ZN(\EXU/CSRControl/_1018_ ) );
AOI21_X1 \EXU/CSRControl/_1876_ ( .A(\EXU/CSRControl/_0978_ ), .B1(\EXU/CSRControl/_1017_ ), .B2(\EXU/CSRControl/_1018_ ), .ZN(\EXU/CSRControl/_1019_ ) );
AOI21_X1 \EXU/CSRControl/_1877_ ( .A(\EXU/CSRControl/_1019_ ), .B1(\EXU/CSRControl/_0205_ ), .B2(\EXU/CSRControl/_0946_ ), .ZN(\EXU/CSRControl/_1020_ ) );
AOI211_X2 \EXU/CSRControl/_1878_ ( .A(\EXU/CSRControl/_0936_ ), .B(\EXU/CSRControl/_1012_ ), .C1(\EXU/CSRControl/_1020_ ), .C2(\EXU/CSRControl/_0935_ ), .ZN(\EXU/CSRControl/_0316_ ) );
BUF_X4 \EXU/CSRControl/_1879_ ( .A(\EXU/CSRControl/_0800_ ), .Z(\EXU/CSRControl/_1021_ ) );
NOR4_X1 \EXU/CSRControl/_1880_ ( .A1(\EXU/CSRControl/_1021_ ), .A2(fanout_net_18 ), .A3(fanout_net_17 ), .A4(\EXU/CSRControl/_0174_ ), .ZN(\EXU/CSRControl/_1022_ ) );
NAND3_X1 \EXU/CSRControl/_1881_ ( .A1(\EXU/CSRControl/_0813_ ), .A2(\EXU/CSRControl/_0174_ ), .A3(\EXU/CSRControl/_0822_ ), .ZN(\EXU/CSRControl/_1023_ ) );
NAND3_X1 \EXU/CSRControl/_1882_ ( .A1(\EXU/CSRControl/_0821_ ), .A2(\EXU/CSRControl/_0238_ ), .A3(\EXU/CSRControl/_0846_ ), .ZN(\EXU/CSRControl/_1024_ ) );
NAND4_X1 \EXU/CSRControl/_1883_ ( .A1(\EXU/CSRControl/_0903_ ), .A2(\EXU/CSRControl/_0829_ ), .A3(\EXU/CSRControl/_0206_ ), .A4(\EXU/CSRControl/_0830_ ), .ZN(\EXU/CSRControl/_1025_ ) );
AND3_X1 \EXU/CSRControl/_1884_ ( .A1(\EXU/CSRControl/_1023_ ), .A2(\EXU/CSRControl/_1024_ ), .A3(\EXU/CSRControl/_1025_ ), .ZN(\EXU/CSRControl/_1026_ ) );
NAND3_X1 \EXU/CSRControl/_1885_ ( .A1(\EXU/CSRControl/_0942_ ), .A2(\EXU/CSRControl/_0142_ ), .A3(\EXU/CSRControl/_0943_ ), .ZN(\EXU/CSRControl/_1027_ ) );
AOI21_X1 \EXU/CSRControl/_1886_ ( .A(\EXU/CSRControl/_0978_ ), .B1(\EXU/CSRControl/_1026_ ), .B2(\EXU/CSRControl/_1027_ ), .ZN(\EXU/CSRControl/_1028_ ) );
AOI21_X1 \EXU/CSRControl/_1887_ ( .A(\EXU/CSRControl/_1028_ ), .B1(\EXU/CSRControl/_0206_ ), .B2(\EXU/CSRControl/_0946_ ), .ZN(\EXU/CSRControl/_1029_ ) );
BUF_X4 \EXU/CSRControl/_1888_ ( .A(\EXU/CSRControl/_0842_ ), .Z(\EXU/CSRControl/_1030_ ) );
AOI211_X2 \EXU/CSRControl/_1889_ ( .A(\EXU/CSRControl/_0936_ ), .B(\EXU/CSRControl/_1022_ ), .C1(\EXU/CSRControl/_1029_ ), .C2(\EXU/CSRControl/_1030_ ), .ZN(\EXU/CSRControl/_0317_ ) );
BUF_X4 \EXU/CSRControl/_1890_ ( .A(\EXU/CSRControl/_0797_ ), .Z(\EXU/CSRControl/_1031_ ) );
NOR4_X1 \EXU/CSRControl/_1891_ ( .A1(\EXU/CSRControl/_1021_ ), .A2(fanout_net_18 ), .A3(fanout_net_17 ), .A4(\EXU/CSRControl/_0176_ ), .ZN(\EXU/CSRControl/_1032_ ) );
NAND3_X1 \EXU/CSRControl/_1892_ ( .A1(\EXU/CSRControl/_0957_ ), .A2(\EXU/CSRControl/_0176_ ), .A3(\EXU/CSRControl/_0958_ ), .ZN(\EXU/CSRControl/_1033_ ) );
NAND3_X1 \EXU/CSRControl/_1893_ ( .A1(\EXU/CSRControl/_0969_ ), .A2(\EXU/CSRControl/_0240_ ), .A3(\EXU/CSRControl/_0960_ ), .ZN(\EXU/CSRControl/_1034_ ) );
NAND4_X1 \EXU/CSRControl/_1894_ ( .A1(\EXU/CSRControl/_0981_ ), .A2(\EXU/CSRControl/_0971_ ), .A3(\EXU/CSRControl/_0208_ ), .A4(\EXU/CSRControl/_0982_ ), .ZN(\EXU/CSRControl/_1035_ ) );
AND4_X1 \EXU/CSRControl/_1895_ ( .A1(\EXU/CSRControl/_0866_ ), .A2(\EXU/CSRControl/_1033_ ), .A3(\EXU/CSRControl/_1034_ ), .A4(\EXU/CSRControl/_1035_ ), .ZN(\EXU/CSRControl/_1036_ ) );
BUF_X4 \EXU/CSRControl/_1896_ ( .A(\EXU/CSRControl/_0833_ ), .Z(\EXU/CSRControl/_1037_ ) );
BUF_X4 \EXU/CSRControl/_1897_ ( .A(\EXU/CSRControl/_0816_ ), .Z(\EXU/CSRControl/_1038_ ) );
NAND3_X1 \EXU/CSRControl/_1898_ ( .A1(\EXU/CSRControl/_1037_ ), .A2(\EXU/CSRControl/_0144_ ), .A3(\EXU/CSRControl/_1038_ ), .ZN(\EXU/CSRControl/_1039_ ) );
AOI21_X1 \EXU/CSRControl/_1899_ ( .A(\EXU/CSRControl/_0978_ ), .B1(\EXU/CSRControl/_1036_ ), .B2(\EXU/CSRControl/_1039_ ), .ZN(\EXU/CSRControl/_1040_ ) );
BUF_X4 \EXU/CSRControl/_1900_ ( .A(\EXU/CSRControl/_0805_ ), .Z(\EXU/CSRControl/_1041_ ) );
AOI21_X1 \EXU/CSRControl/_1901_ ( .A(\EXU/CSRControl/_1040_ ), .B1(\EXU/CSRControl/_0208_ ), .B2(\EXU/CSRControl/_1041_ ), .ZN(\EXU/CSRControl/_1042_ ) );
AOI211_X2 \EXU/CSRControl/_1902_ ( .A(\EXU/CSRControl/_1031_ ), .B(\EXU/CSRControl/_1032_ ), .C1(\EXU/CSRControl/_1042_ ), .C2(\EXU/CSRControl/_1030_ ), .ZN(\EXU/CSRControl/_0319_ ) );
NOR4_X1 \EXU/CSRControl/_1903_ ( .A1(\EXU/CSRControl/_1021_ ), .A2(fanout_net_18 ), .A3(fanout_net_17 ), .A4(\EXU/CSRControl/_0177_ ), .ZN(\EXU/CSRControl/_1043_ ) );
NAND3_X1 \EXU/CSRControl/_1904_ ( .A1(\EXU/CSRControl/_0957_ ), .A2(\EXU/CSRControl/_0177_ ), .A3(\EXU/CSRControl/_0958_ ), .ZN(\EXU/CSRControl/_1044_ ) );
NAND3_X1 \EXU/CSRControl/_1905_ ( .A1(\EXU/CSRControl/_0969_ ), .A2(\EXU/CSRControl/_0241_ ), .A3(\EXU/CSRControl/_0960_ ), .ZN(\EXU/CSRControl/_1045_ ) );
NAND4_X1 \EXU/CSRControl/_1906_ ( .A1(\EXU/CSRControl/_0981_ ), .A2(\EXU/CSRControl/_0971_ ), .A3(\EXU/CSRControl/_0209_ ), .A4(\EXU/CSRControl/_0982_ ), .ZN(\EXU/CSRControl/_1046_ ) );
AND4_X1 \EXU/CSRControl/_1907_ ( .A1(\EXU/CSRControl/_0866_ ), .A2(\EXU/CSRControl/_1044_ ), .A3(\EXU/CSRControl/_1045_ ), .A4(\EXU/CSRControl/_1046_ ), .ZN(\EXU/CSRControl/_1047_ ) );
NAND3_X1 \EXU/CSRControl/_1908_ ( .A1(\EXU/CSRControl/_1037_ ), .A2(\EXU/CSRControl/_0145_ ), .A3(\EXU/CSRControl/_1038_ ), .ZN(\EXU/CSRControl/_1048_ ) );
AOI21_X1 \EXU/CSRControl/_1909_ ( .A(\EXU/CSRControl/_0978_ ), .B1(\EXU/CSRControl/_1047_ ), .B2(\EXU/CSRControl/_1048_ ), .ZN(\EXU/CSRControl/_1049_ ) );
AOI21_X1 \EXU/CSRControl/_1910_ ( .A(\EXU/CSRControl/_1049_ ), .B1(\EXU/CSRControl/_0209_ ), .B2(\EXU/CSRControl/_1041_ ), .ZN(\EXU/CSRControl/_1050_ ) );
AOI211_X2 \EXU/CSRControl/_1911_ ( .A(\EXU/CSRControl/_1031_ ), .B(\EXU/CSRControl/_1043_ ), .C1(\EXU/CSRControl/_1050_ ), .C2(\EXU/CSRControl/_1030_ ), .ZN(\EXU/CSRControl/_0320_ ) );
NOR4_X1 \EXU/CSRControl/_1912_ ( .A1(\EXU/CSRControl/_1021_ ), .A2(fanout_net_18 ), .A3(fanout_net_17 ), .A4(\EXU/CSRControl/_0178_ ), .ZN(\EXU/CSRControl/_1051_ ) );
NAND3_X1 \EXU/CSRControl/_1913_ ( .A1(\EXU/CSRControl/_0957_ ), .A2(\EXU/CSRControl/_0178_ ), .A3(\EXU/CSRControl/_0958_ ), .ZN(\EXU/CSRControl/_1052_ ) );
NAND3_X1 \EXU/CSRControl/_1914_ ( .A1(\EXU/CSRControl/_0969_ ), .A2(\EXU/CSRControl/_0242_ ), .A3(\EXU/CSRControl/_0960_ ), .ZN(\EXU/CSRControl/_1053_ ) );
NAND4_X1 \EXU/CSRControl/_1915_ ( .A1(\EXU/CSRControl/_0981_ ), .A2(\EXU/CSRControl/_0971_ ), .A3(\EXU/CSRControl/_0210_ ), .A4(\EXU/CSRControl/_0982_ ), .ZN(\EXU/CSRControl/_1054_ ) );
AND4_X1 \EXU/CSRControl/_1916_ ( .A1(\EXU/CSRControl/_0866_ ), .A2(\EXU/CSRControl/_1052_ ), .A3(\EXU/CSRControl/_1053_ ), .A4(\EXU/CSRControl/_1054_ ), .ZN(\EXU/CSRControl/_1055_ ) );
NAND3_X1 \EXU/CSRControl/_1917_ ( .A1(\EXU/CSRControl/_1037_ ), .A2(\EXU/CSRControl/_0146_ ), .A3(\EXU/CSRControl/_1038_ ), .ZN(\EXU/CSRControl/_1056_ ) );
AOI21_X1 \EXU/CSRControl/_1918_ ( .A(\EXU/CSRControl/_0978_ ), .B1(\EXU/CSRControl/_1055_ ), .B2(\EXU/CSRControl/_1056_ ), .ZN(\EXU/CSRControl/_1057_ ) );
AOI21_X1 \EXU/CSRControl/_1919_ ( .A(\EXU/CSRControl/_1057_ ), .B1(\EXU/CSRControl/_0210_ ), .B2(\EXU/CSRControl/_1041_ ), .ZN(\EXU/CSRControl/_1058_ ) );
AOI211_X2 \EXU/CSRControl/_1920_ ( .A(\EXU/CSRControl/_1031_ ), .B(\EXU/CSRControl/_1051_ ), .C1(\EXU/CSRControl/_1058_ ), .C2(\EXU/CSRControl/_1030_ ), .ZN(\EXU/CSRControl/_0321_ ) );
NOR4_X1 \EXU/CSRControl/_1921_ ( .A1(\EXU/CSRControl/_1021_ ), .A2(fanout_net_18 ), .A3(fanout_net_17 ), .A4(\EXU/CSRControl/_0179_ ), .ZN(\EXU/CSRControl/_1059_ ) );
NAND3_X1 \EXU/CSRControl/_1922_ ( .A1(\EXU/CSRControl/_0813_ ), .A2(\EXU/CSRControl/_0179_ ), .A3(\EXU/CSRControl/_0822_ ), .ZN(\EXU/CSRControl/_1060_ ) );
NAND3_X1 \EXU/CSRControl/_1923_ ( .A1(\EXU/CSRControl/_0821_ ), .A2(\EXU/CSRControl/_0243_ ), .A3(\EXU/CSRControl/_0846_ ), .ZN(\EXU/CSRControl/_1061_ ) );
NAND4_X1 \EXU/CSRControl/_1924_ ( .A1(\EXU/CSRControl/_0903_ ), .A2(\EXU/CSRControl/_0829_ ), .A3(\EXU/CSRControl/_0211_ ), .A4(\EXU/CSRControl/_0872_ ), .ZN(\EXU/CSRControl/_1062_ ) );
AND3_X1 \EXU/CSRControl/_1925_ ( .A1(\EXU/CSRControl/_1060_ ), .A2(\EXU/CSRControl/_1061_ ), .A3(\EXU/CSRControl/_1062_ ), .ZN(\EXU/CSRControl/_1063_ ) );
NAND3_X1 \EXU/CSRControl/_1926_ ( .A1(\EXU/CSRControl/_1037_ ), .A2(\EXU/CSRControl/_0147_ ), .A3(\EXU/CSRControl/_1038_ ), .ZN(\EXU/CSRControl/_1064_ ) );
AOI21_X1 \EXU/CSRControl/_1927_ ( .A(\EXU/CSRControl/_0978_ ), .B1(\EXU/CSRControl/_1063_ ), .B2(\EXU/CSRControl/_1064_ ), .ZN(\EXU/CSRControl/_1065_ ) );
AOI21_X1 \EXU/CSRControl/_1928_ ( .A(\EXU/CSRControl/_1065_ ), .B1(\EXU/CSRControl/_0211_ ), .B2(\EXU/CSRControl/_1041_ ), .ZN(\EXU/CSRControl/_1066_ ) );
AOI211_X2 \EXU/CSRControl/_1929_ ( .A(\EXU/CSRControl/_1031_ ), .B(\EXU/CSRControl/_1059_ ), .C1(\EXU/CSRControl/_1066_ ), .C2(\EXU/CSRControl/_1030_ ), .ZN(\EXU/CSRControl/_0322_ ) );
NOR4_X1 \EXU/CSRControl/_1930_ ( .A1(\EXU/CSRControl/_1021_ ), .A2(fanout_net_18 ), .A3(fanout_net_17 ), .A4(\EXU/CSRControl/_0180_ ), .ZN(\EXU/CSRControl/_1067_ ) );
NAND3_X1 \EXU/CSRControl/_1931_ ( .A1(\EXU/CSRControl/_0957_ ), .A2(\EXU/CSRControl/_0180_ ), .A3(\EXU/CSRControl/_0958_ ), .ZN(\EXU/CSRControl/_1068_ ) );
NAND3_X1 \EXU/CSRControl/_1932_ ( .A1(\EXU/CSRControl/_0969_ ), .A2(\EXU/CSRControl/_0244_ ), .A3(\EXU/CSRControl/_0960_ ), .ZN(\EXU/CSRControl/_1069_ ) );
NAND4_X1 \EXU/CSRControl/_1933_ ( .A1(\EXU/CSRControl/_0981_ ), .A2(\EXU/CSRControl/_0971_ ), .A3(\EXU/CSRControl/_0212_ ), .A4(\EXU/CSRControl/_0982_ ), .ZN(\EXU/CSRControl/_1070_ ) );
AND4_X1 \EXU/CSRControl/_1934_ ( .A1(\EXU/CSRControl/_0866_ ), .A2(\EXU/CSRControl/_1068_ ), .A3(\EXU/CSRControl/_1069_ ), .A4(\EXU/CSRControl/_1070_ ), .ZN(\EXU/CSRControl/_1071_ ) );
NAND3_X1 \EXU/CSRControl/_1935_ ( .A1(\EXU/CSRControl/_1037_ ), .A2(\EXU/CSRControl/_0148_ ), .A3(\EXU/CSRControl/_1038_ ), .ZN(\EXU/CSRControl/_1072_ ) );
AOI21_X1 \EXU/CSRControl/_1936_ ( .A(\EXU/CSRControl/_0883_ ), .B1(\EXU/CSRControl/_1071_ ), .B2(\EXU/CSRControl/_1072_ ), .ZN(\EXU/CSRControl/_1073_ ) );
AOI21_X1 \EXU/CSRControl/_1937_ ( .A(\EXU/CSRControl/_1073_ ), .B1(\EXU/CSRControl/_0212_ ), .B2(\EXU/CSRControl/_1041_ ), .ZN(\EXU/CSRControl/_1074_ ) );
AOI211_X2 \EXU/CSRControl/_1938_ ( .A(\EXU/CSRControl/_1031_ ), .B(\EXU/CSRControl/_1067_ ), .C1(\EXU/CSRControl/_1074_ ), .C2(\EXU/CSRControl/_1030_ ), .ZN(\EXU/CSRControl/_0323_ ) );
NOR4_X1 \EXU/CSRControl/_1939_ ( .A1(\EXU/CSRControl/_1021_ ), .A2(fanout_net_18 ), .A3(fanout_net_17 ), .A4(\EXU/CSRControl/_0181_ ), .ZN(\EXU/CSRControl/_1075_ ) );
NAND3_X1 \EXU/CSRControl/_1940_ ( .A1(\EXU/CSRControl/_0813_ ), .A2(\EXU/CSRControl/_0181_ ), .A3(\EXU/CSRControl/_0822_ ), .ZN(\EXU/CSRControl/_1076_ ) );
NAND3_X1 \EXU/CSRControl/_1941_ ( .A1(\EXU/CSRControl/_0821_ ), .A2(\EXU/CSRControl/_0245_ ), .A3(\EXU/CSRControl/_0846_ ), .ZN(\EXU/CSRControl/_1077_ ) );
NAND4_X1 \EXU/CSRControl/_1942_ ( .A1(\EXU/CSRControl/_0903_ ), .A2(\EXU/CSRControl/_0875_ ), .A3(\EXU/CSRControl/_0213_ ), .A4(\EXU/CSRControl/_0872_ ), .ZN(\EXU/CSRControl/_1078_ ) );
AND3_X1 \EXU/CSRControl/_1943_ ( .A1(\EXU/CSRControl/_1076_ ), .A2(\EXU/CSRControl/_1077_ ), .A3(\EXU/CSRControl/_1078_ ), .ZN(\EXU/CSRControl/_1079_ ) );
NAND3_X1 \EXU/CSRControl/_1944_ ( .A1(\EXU/CSRControl/_1037_ ), .A2(\EXU/CSRControl/_0149_ ), .A3(\EXU/CSRControl/_1038_ ), .ZN(\EXU/CSRControl/_1080_ ) );
AOI21_X1 \EXU/CSRControl/_1945_ ( .A(\EXU/CSRControl/_0883_ ), .B1(\EXU/CSRControl/_1079_ ), .B2(\EXU/CSRControl/_1080_ ), .ZN(\EXU/CSRControl/_1081_ ) );
AOI21_X1 \EXU/CSRControl/_1946_ ( .A(\EXU/CSRControl/_1081_ ), .B1(\EXU/CSRControl/_0213_ ), .B2(\EXU/CSRControl/_1041_ ), .ZN(\EXU/CSRControl/_1082_ ) );
AOI211_X2 \EXU/CSRControl/_1947_ ( .A(\EXU/CSRControl/_1031_ ), .B(\EXU/CSRControl/_1075_ ), .C1(\EXU/CSRControl/_1082_ ), .C2(\EXU/CSRControl/_1030_ ), .ZN(\EXU/CSRControl/_0324_ ) );
NOR4_X1 \EXU/CSRControl/_1948_ ( .A1(\EXU/CSRControl/_1021_ ), .A2(fanout_net_18 ), .A3(fanout_net_17 ), .A4(\EXU/CSRControl/_0182_ ), .ZN(\EXU/CSRControl/_1083_ ) );
NAND3_X1 \EXU/CSRControl/_1949_ ( .A1(\EXU/CSRControl/_0868_ ), .A2(\EXU/CSRControl/_0182_ ), .A3(\EXU/CSRControl/_0822_ ), .ZN(\EXU/CSRControl/_1084_ ) );
NAND3_X1 \EXU/CSRControl/_1950_ ( .A1(\EXU/CSRControl/_0871_ ), .A2(\EXU/CSRControl/_0246_ ), .A3(\EXU/CSRControl/_0846_ ), .ZN(\EXU/CSRControl/_1085_ ) );
NAND4_X1 \EXU/CSRControl/_1951_ ( .A1(\EXU/CSRControl/_0903_ ), .A2(\EXU/CSRControl/_0875_ ), .A3(\EXU/CSRControl/_0214_ ), .A4(\EXU/CSRControl/_0872_ ), .ZN(\EXU/CSRControl/_1086_ ) );
AND3_X1 \EXU/CSRControl/_1952_ ( .A1(\EXU/CSRControl/_1084_ ), .A2(\EXU/CSRControl/_1085_ ), .A3(\EXU/CSRControl/_1086_ ), .ZN(\EXU/CSRControl/_1087_ ) );
NAND3_X1 \EXU/CSRControl/_1953_ ( .A1(\EXU/CSRControl/_1037_ ), .A2(\EXU/CSRControl/_0150_ ), .A3(\EXU/CSRControl/_1038_ ), .ZN(\EXU/CSRControl/_1088_ ) );
AOI21_X1 \EXU/CSRControl/_1954_ ( .A(\EXU/CSRControl/_0883_ ), .B1(\EXU/CSRControl/_1087_ ), .B2(\EXU/CSRControl/_1088_ ), .ZN(\EXU/CSRControl/_1089_ ) );
AOI21_X1 \EXU/CSRControl/_1955_ ( .A(\EXU/CSRControl/_1089_ ), .B1(\EXU/CSRControl/_0214_ ), .B2(\EXU/CSRControl/_1041_ ), .ZN(\EXU/CSRControl/_1090_ ) );
AOI211_X2 \EXU/CSRControl/_1956_ ( .A(\EXU/CSRControl/_1031_ ), .B(\EXU/CSRControl/_1083_ ), .C1(\EXU/CSRControl/_1090_ ), .C2(\EXU/CSRControl/_1030_ ), .ZN(\EXU/CSRControl/_0325_ ) );
NOR4_X1 \EXU/CSRControl/_1957_ ( .A1(\EXU/CSRControl/_1021_ ), .A2(fanout_net_18 ), .A3(fanout_net_17 ), .A4(\EXU/CSRControl/_0183_ ), .ZN(\EXU/CSRControl/_1091_ ) );
NAND3_X1 \EXU/CSRControl/_1958_ ( .A1(\EXU/CSRControl/_0957_ ), .A2(\EXU/CSRControl/_0183_ ), .A3(\EXU/CSRControl/_0958_ ), .ZN(\EXU/CSRControl/_1092_ ) );
NAND3_X1 \EXU/CSRControl/_1959_ ( .A1(\EXU/CSRControl/_0969_ ), .A2(\EXU/CSRControl/_0247_ ), .A3(\EXU/CSRControl/_0960_ ), .ZN(\EXU/CSRControl/_1093_ ) );
NAND4_X1 \EXU/CSRControl/_1960_ ( .A1(\EXU/CSRControl/_0981_ ), .A2(\EXU/CSRControl/_0971_ ), .A3(\EXU/CSRControl/_0215_ ), .A4(\EXU/CSRControl/_0982_ ), .ZN(\EXU/CSRControl/_1094_ ) );
AND4_X1 \EXU/CSRControl/_1961_ ( .A1(\EXU/CSRControl/_0866_ ), .A2(\EXU/CSRControl/_1092_ ), .A3(\EXU/CSRControl/_1093_ ), .A4(\EXU/CSRControl/_1094_ ), .ZN(\EXU/CSRControl/_1095_ ) );
NAND3_X1 \EXU/CSRControl/_1962_ ( .A1(\EXU/CSRControl/_1037_ ), .A2(\EXU/CSRControl/_0151_ ), .A3(\EXU/CSRControl/_1038_ ), .ZN(\EXU/CSRControl/_1096_ ) );
AOI21_X1 \EXU/CSRControl/_1963_ ( .A(\EXU/CSRControl/_0883_ ), .B1(\EXU/CSRControl/_1095_ ), .B2(\EXU/CSRControl/_1096_ ), .ZN(\EXU/CSRControl/_1097_ ) );
AOI21_X1 \EXU/CSRControl/_1964_ ( .A(\EXU/CSRControl/_1097_ ), .B1(\EXU/CSRControl/_0215_ ), .B2(\EXU/CSRControl/_1041_ ), .ZN(\EXU/CSRControl/_1098_ ) );
AOI211_X2 \EXU/CSRControl/_1965_ ( .A(\EXU/CSRControl/_1031_ ), .B(\EXU/CSRControl/_1091_ ), .C1(\EXU/CSRControl/_1098_ ), .C2(\EXU/CSRControl/_1030_ ), .ZN(\EXU/CSRControl/_0326_ ) );
NOR4_X1 \EXU/CSRControl/_1966_ ( .A1(\EXU/CSRControl/_1021_ ), .A2(\EXU/CSRControl/_0273_ ), .A3(\EXU/CSRControl/_0272_ ), .A4(\EXU/CSRControl/_0184_ ), .ZN(\EXU/CSRControl/_1099_ ) );
NAND3_X1 \EXU/CSRControl/_1967_ ( .A1(\EXU/CSRControl/_0812_ ), .A2(\EXU/CSRControl/_0184_ ), .A3(\EXU/CSRControl/_0830_ ), .ZN(\EXU/CSRControl/_1100_ ) );
NAND3_X1 \EXU/CSRControl/_1968_ ( .A1(\EXU/CSRControl/_0969_ ), .A2(\EXU/CSRControl/_0248_ ), .A3(\EXU/CSRControl/_0876_ ), .ZN(\EXU/CSRControl/_1101_ ) );
NAND4_X1 \EXU/CSRControl/_1969_ ( .A1(\EXU/CSRControl/_0981_ ), .A2(\EXU/CSRControl/_0971_ ), .A3(\EXU/CSRControl/_0216_ ), .A4(\EXU/CSRControl/_0982_ ), .ZN(\EXU/CSRControl/_1102_ ) );
AND4_X1 \EXU/CSRControl/_1970_ ( .A1(\EXU/CSRControl/_0866_ ), .A2(\EXU/CSRControl/_1100_ ), .A3(\EXU/CSRControl/_1101_ ), .A4(\EXU/CSRControl/_1102_ ), .ZN(\EXU/CSRControl/_1103_ ) );
NAND3_X1 \EXU/CSRControl/_1971_ ( .A1(\EXU/CSRControl/_1037_ ), .A2(\EXU/CSRControl/_0152_ ), .A3(\EXU/CSRControl/_1038_ ), .ZN(\EXU/CSRControl/_1104_ ) );
AOI21_X1 \EXU/CSRControl/_1972_ ( .A(\EXU/CSRControl/_0883_ ), .B1(\EXU/CSRControl/_1103_ ), .B2(\EXU/CSRControl/_1104_ ), .ZN(\EXU/CSRControl/_1105_ ) );
AOI21_X1 \EXU/CSRControl/_1973_ ( .A(\EXU/CSRControl/_1105_ ), .B1(\EXU/CSRControl/_0216_ ), .B2(\EXU/CSRControl/_1041_ ), .ZN(\EXU/CSRControl/_1106_ ) );
AOI211_X2 \EXU/CSRControl/_1974_ ( .A(\EXU/CSRControl/_1031_ ), .B(\EXU/CSRControl/_1099_ ), .C1(\EXU/CSRControl/_1106_ ), .C2(\EXU/CSRControl/_1030_ ), .ZN(\EXU/CSRControl/_0327_ ) );
NOR4_X1 \EXU/CSRControl/_1975_ ( .A1(\EXU/CSRControl/_0800_ ), .A2(\EXU/CSRControl/_0273_ ), .A3(\EXU/CSRControl/_0272_ ), .A4(\EXU/CSRControl/_0185_ ), .ZN(\EXU/CSRControl/_1107_ ) );
NAND3_X1 \EXU/CSRControl/_1976_ ( .A1(\EXU/CSRControl/_0812_ ), .A2(\EXU/CSRControl/_0185_ ), .A3(\EXU/CSRControl/_0830_ ), .ZN(\EXU/CSRControl/_1108_ ) );
NAND3_X1 \EXU/CSRControl/_1977_ ( .A1(\EXU/CSRControl/_0820_ ), .A2(\EXU/CSRControl/_0249_ ), .A3(\EXU/CSRControl/_0876_ ), .ZN(\EXU/CSRControl/_1109_ ) );
NAND4_X1 \EXU/CSRControl/_1978_ ( .A1(\EXU/CSRControl/_0981_ ), .A2(\EXU/CSRControl/_0828_ ), .A3(\EXU/CSRControl/_0217_ ), .A4(\EXU/CSRControl/_0982_ ), .ZN(\EXU/CSRControl/_1110_ ) );
AND4_X1 \EXU/CSRControl/_1979_ ( .A1(\EXU/CSRControl/_0866_ ), .A2(\EXU/CSRControl/_1108_ ), .A3(\EXU/CSRControl/_1109_ ), .A4(\EXU/CSRControl/_1110_ ), .ZN(\EXU/CSRControl/_1111_ ) );
NAND3_X1 \EXU/CSRControl/_1980_ ( .A1(\EXU/CSRControl/_1037_ ), .A2(\EXU/CSRControl/_0153_ ), .A3(\EXU/CSRControl/_1038_ ), .ZN(\EXU/CSRControl/_1112_ ) );
AOI21_X1 \EXU/CSRControl/_1981_ ( .A(\EXU/CSRControl/_0883_ ), .B1(\EXU/CSRControl/_1111_ ), .B2(\EXU/CSRControl/_1112_ ), .ZN(\EXU/CSRControl/_1113_ ) );
AOI21_X1 \EXU/CSRControl/_1982_ ( .A(\EXU/CSRControl/_1113_ ), .B1(\EXU/CSRControl/_0217_ ), .B2(\EXU/CSRControl/_1041_ ), .ZN(\EXU/CSRControl/_1114_ ) );
AOI211_X2 \EXU/CSRControl/_1983_ ( .A(\EXU/CSRControl/_1031_ ), .B(\EXU/CSRControl/_1107_ ), .C1(\EXU/CSRControl/_1114_ ), .C2(\EXU/CSRControl/_0842_ ), .ZN(\EXU/CSRControl/_0328_ ) );
NOR4_X1 \EXU/CSRControl/_1984_ ( .A1(\EXU/CSRControl/_0800_ ), .A2(\EXU/CSRControl/_0273_ ), .A3(\EXU/CSRControl/_0272_ ), .A4(\EXU/CSRControl/_0187_ ), .ZN(\EXU/CSRControl/_1115_ ) );
AND3_X1 \EXU/CSRControl/_1985_ ( .A1(\EXU/CSRControl/_0868_ ), .A2(\EXU/CSRControl/_0187_ ), .A3(\EXU/CSRControl/_0869_ ), .ZN(\EXU/CSRControl/_1116_ ) );
BUF_X4 \EXU/CSRControl/_1986_ ( .A(\EXU/CSRControl/_0826_ ), .Z(\EXU/CSRControl/_1117_ ) );
NAND4_X1 \EXU/CSRControl/_1987_ ( .A1(\EXU/CSRControl/_1117_ ), .A2(\EXU/CSRControl/_0828_ ), .A3(\EXU/CSRControl/_0219_ ), .A4(\EXU/CSRControl/_0815_ ), .ZN(\EXU/CSRControl/_1118_ ) );
NAND3_X1 \EXU/CSRControl/_1988_ ( .A1(\EXU/CSRControl/_0820_ ), .A2(\EXU/CSRControl/_0251_ ), .A3(\EXU/CSRControl/_0876_ ), .ZN(\EXU/CSRControl/_1119_ ) );
NAND2_X1 \EXU/CSRControl/_1989_ ( .A1(\EXU/CSRControl/_1118_ ), .A2(\EXU/CSRControl/_1119_ ), .ZN(\EXU/CSRControl/_1120_ ) );
NOR3_X1 \EXU/CSRControl/_1990_ ( .A1(\EXU/CSRControl/_1116_ ), .A2(\EXU/CSRControl/_0865_ ), .A3(\EXU/CSRControl/_1120_ ), .ZN(\EXU/CSRControl/_1121_ ) );
NAND3_X1 \EXU/CSRControl/_1991_ ( .A1(\EXU/CSRControl/_0833_ ), .A2(\EXU/CSRControl/_0155_ ), .A3(\EXU/CSRControl/_0816_ ), .ZN(\EXU/CSRControl/_1122_ ) );
AOI21_X1 \EXU/CSRControl/_1992_ ( .A(\EXU/CSRControl/_0883_ ), .B1(\EXU/CSRControl/_1121_ ), .B2(\EXU/CSRControl/_1122_ ), .ZN(\EXU/CSRControl/_1123_ ) );
AOI21_X1 \EXU/CSRControl/_1993_ ( .A(\EXU/CSRControl/_1123_ ), .B1(\EXU/CSRControl/_0219_ ), .B2(\EXU/CSRControl/_0805_ ), .ZN(\EXU/CSRControl/_1124_ ) );
AOI211_X2 \EXU/CSRControl/_1994_ ( .A(\EXU/CSRControl/_0797_ ), .B(\EXU/CSRControl/_1115_ ), .C1(\EXU/CSRControl/_1124_ ), .C2(\EXU/CSRControl/_0842_ ), .ZN(\EXU/CSRControl/_0330_ ) );
NOR4_X1 \EXU/CSRControl/_1995_ ( .A1(\EXU/CSRControl/_0800_ ), .A2(\EXU/CSRControl/_0273_ ), .A3(\EXU/CSRControl/_0272_ ), .A4(\EXU/CSRControl/_0188_ ), .ZN(\EXU/CSRControl/_1125_ ) );
NAND3_X1 \EXU/CSRControl/_1996_ ( .A1(\EXU/CSRControl/_0868_ ), .A2(\EXU/CSRControl/_0188_ ), .A3(\EXU/CSRControl/_0822_ ), .ZN(\EXU/CSRControl/_1126_ ) );
NAND3_X1 \EXU/CSRControl/_1997_ ( .A1(\EXU/CSRControl/_0871_ ), .A2(\EXU/CSRControl/_0252_ ), .A3(\EXU/CSRControl/_0869_ ), .ZN(\EXU/CSRControl/_1127_ ) );
NAND4_X1 \EXU/CSRControl/_1998_ ( .A1(\EXU/CSRControl/_0903_ ), .A2(\EXU/CSRControl/_0875_ ), .A3(\EXU/CSRControl/_0220_ ), .A4(\EXU/CSRControl/_0872_ ), .ZN(\EXU/CSRControl/_1128_ ) );
AND3_X1 \EXU/CSRControl/_1999_ ( .A1(\EXU/CSRControl/_1126_ ), .A2(\EXU/CSRControl/_1127_ ), .A3(\EXU/CSRControl/_1128_ ), .ZN(\EXU/CSRControl/_1129_ ) );
NAND3_X1 \EXU/CSRControl/_2000_ ( .A1(\EXU/CSRControl/_0833_ ), .A2(\EXU/CSRControl/_0156_ ), .A3(\EXU/CSRControl/_0816_ ), .ZN(\EXU/CSRControl/_1130_ ) );
AOI21_X1 \EXU/CSRControl/_2001_ ( .A(\EXU/CSRControl/_0883_ ), .B1(\EXU/CSRControl/_1129_ ), .B2(\EXU/CSRControl/_1130_ ), .ZN(\EXU/CSRControl/_1131_ ) );
AOI21_X1 \EXU/CSRControl/_2002_ ( .A(\EXU/CSRControl/_1131_ ), .B1(\EXU/CSRControl/_0220_ ), .B2(\EXU/CSRControl/_0805_ ), .ZN(\EXU/CSRControl/_1132_ ) );
AOI211_X4 \EXU/CSRControl/_2003_ ( .A(\EXU/CSRControl/_0797_ ), .B(\EXU/CSRControl/_1125_ ), .C1(\EXU/CSRControl/_1132_ ), .C2(\EXU/CSRControl/_0842_ ), .ZN(\EXU/CSRControl/_0331_ ) );
AND2_X1 \EXU/CSRControl/_2004_ ( .A1(\EXU/CSRControl/_0796_ ), .A2(\EXU/CSRControl/_0272_ ), .ZN(\EXU/CSRControl/_1133_ ) );
INV_X1 \EXU/CSRControl/_2005_ ( .A(\EXU/CSRControl/_1133_ ), .ZN(\EXU/CSRControl/_1134_ ) );
OR2_X2 \EXU/CSRControl/_2006_ ( .A1(\EXU/CSRControl/_1134_ ), .A2(\EXU/CSRControl/_0273_ ), .ZN(\EXU/CSRControl/_1135_ ) );
NAND3_X1 \EXU/CSRControl/_2007_ ( .A1(\EXU/CSRControl/_0796_ ), .A2(\EXU/CSRControl/_0272_ ), .A3(\EXU/CSRControl/_0300_ ), .ZN(\EXU/CSRControl/_1136_ ) );
INV_X8 \EXU/CSRControl/_2008_ ( .A(\EXU/CSRControl/_0809_ ), .ZN(\EXU/CSRControl/_1137_ ) );
NAND3_X4 \EXU/CSRControl/_2009_ ( .A1(\EXU/CSRControl/_0814_ ), .A2(\EXU/CSRControl/_0818_ ), .A3(\EXU/CSRControl/_0819_ ), .ZN(\EXU/CSRControl/_1138_ ) );
NOR2_X4 \EXU/CSRControl/_2010_ ( .A1(\EXU/CSRControl/_1137_ ), .A2(\EXU/CSRControl/_1138_ ), .ZN(\EXU/CSRControl/_1139_ ) );
NAND2_X1 \EXU/CSRControl/_2011_ ( .A1(\EXU/CSRControl/_1139_ ), .A2(\EXU/CSRControl/_0253_ ), .ZN(\EXU/CSRControl/_1140_ ) );
AND3_X4 \EXU/CSRControl/_2012_ ( .A1(\EXU/CSRControl/_0811_ ), .A2(\EXU/CSRControl/_0814_ ), .A3(\EXU/CSRControl/_0818_ ), .ZN(\EXU/CSRControl/_1141_ ) );
NAND3_X1 \EXU/CSRControl/_2013_ ( .A1(\EXU/CSRControl/_1141_ ), .A2(\EXU/CSRControl/_0826_ ), .A3(\EXU/CSRControl/_0221_ ), .ZN(\EXU/CSRControl/_1142_ ) );
AND4_X4 \EXU/CSRControl/_2014_ ( .A1(\EXU/CSRControl/_0263_ ), .A2(\EXU/CSRControl/_0814_ ), .A3(\EXU/CSRControl/_0810_ ), .A4(\EXU/CSRControl/_0818_ ), .ZN(\EXU/CSRControl/_1143_ ) );
NAND3_X1 \EXU/CSRControl/_2015_ ( .A1(\EXU/CSRControl/_1143_ ), .A2(\EXU/CSRControl/_0826_ ), .A3(\EXU/CSRControl/_0157_ ), .ZN(\EXU/CSRControl/_1144_ ) );
NAND3_X2 \EXU/CSRControl/_2016_ ( .A1(\EXU/CSRControl/_1140_ ), .A2(\EXU/CSRControl/_1142_ ), .A3(\EXU/CSRControl/_1144_ ), .ZN(\EXU/CSRControl/_1145_ ) );
NAND4_X2 \EXU/CSRControl/_2017_ ( .A1(\EXU/CSRControl/_0862_ ), .A2(\EXU/CSRControl/_0266_ ), .A3(\EXU/CSRControl/_0262_ ), .A4(\EXU/CSRControl/_0261_ ), .ZN(\EXU/CSRControl/_1146_ ) );
NOR3_X4 \EXU/CSRControl/_2018_ ( .A1(\EXU/CSRControl/_1146_ ), .A2(\EXU/CSRControl/_0269_ ), .A3(\EXU/CSRControl/_0268_ ), .ZN(\EXU/CSRControl/_1147_ ) );
AND2_X4 \EXU/CSRControl/_2019_ ( .A1(\EXU/CSRControl/_1147_ ), .A2(\EXU/CSRControl/_1141_ ), .ZN(\EXU/CSRControl/_1148_ ) );
INV_X8 \EXU/CSRControl/_2020_ ( .A(\EXU/CSRControl/_1148_ ), .ZN(\EXU/CSRControl/_1149_ ) );
AND4_X4 \EXU/CSRControl/_2021_ ( .A1(\EXU/CSRControl/_0806_ ), .A2(\EXU/CSRControl/_0811_ ), .A3(\EXU/CSRControl/_0264_ ), .A4(\EXU/CSRControl/_0814_ ), .ZN(\EXU/CSRControl/_1150_ ) );
NAND3_X4 \EXU/CSRControl/_2022_ ( .A1(\EXU/CSRControl/_1150_ ), .A2(\EXU/CSRControl/_0189_ ), .A3(\EXU/CSRControl/_0809_ ), .ZN(\EXU/CSRControl/_1151_ ) );
NAND2_X4 \EXU/CSRControl/_2023_ ( .A1(\EXU/CSRControl/_1149_ ), .A2(\EXU/CSRControl/_1151_ ), .ZN(\EXU/CSRControl/_1152_ ) );
OAI211_X4 \EXU/CSRControl/_2024_ ( .A(\EXU/CSRControl/_1135_ ), .B(\EXU/CSRControl/_1136_ ), .C1(\EXU/CSRControl/_1145_ ), .C2(\EXU/CSRControl/_1152_ ), .ZN(\EXU/CSRControl/_1153_ ) );
XNOR2_X1 \EXU/CSRControl/_2025_ ( .A(\EXU/CSRControl/_0273_ ), .B(\EXU/CSRControl/_0272_ ), .ZN(\EXU/CSRControl/_1154_ ) );
NOR2_X1 \EXU/CSRControl/_2026_ ( .A1(\EXU/CSRControl/_1154_ ), .A2(\EXU/CSRControl/_0274_ ), .ZN(\EXU/CSRControl/_1155_ ) );
NAND2_X1 \EXU/CSRControl/_2027_ ( .A1(\EXU/CSRControl/_1155_ ), .A2(\EXU/CSRControl/_0300_ ), .ZN(\EXU/CSRControl/_1156_ ) );
AND2_X4 \EXU/CSRControl/_2028_ ( .A1(\EXU/CSRControl/_1153_ ), .A2(\EXU/CSRControl/_1156_ ), .ZN(\EXU/CSRControl/_1157_ ) );
INV_X1 \EXU/CSRControl/_2029_ ( .A(\EXU/CSRControl/_0883_ ), .ZN(\EXU/CSRControl/_1158_ ) );
MUX2_X2 \EXU/CSRControl/_2030_ ( .A(\EXU/CSRControl/_0001_ ), .B(\EXU/CSRControl/_1157_ ), .S(\EXU/CSRControl/_1158_ ), .Z(\EXU/CSRControl/_1159_ ) );
BUF_X2 \EXU/CSRControl/_2031_ ( .A(\EXU/CSRControl/_0841_ ), .Z(\EXU/CSRControl/_1160_ ) );
NOR3_X2 \EXU/CSRControl/_2032_ ( .A1(\EXU/CSRControl/_1137_ ), .A2(\EXU/CSRControl/_1138_ ), .A3(\EXU/CSRControl/_0795_ ), .ZN(\EXU/CSRControl/_1161_ ) );
NOR2_X1 \EXU/CSRControl/_2033_ ( .A1(\EXU/CSRControl/_1161_ ), .A2(\EXU/CSRControl/_0803_ ), .ZN(\EXU/CSRControl/_1162_ ) );
OR3_X4 \EXU/CSRControl/_2034_ ( .A1(\EXU/CSRControl/_1159_ ), .A2(\EXU/CSRControl/_1160_ ), .A3(\EXU/CSRControl/_1162_ ), .ZN(\EXU/CSRControl/_1163_ ) );
NAND2_X1 \EXU/CSRControl/_2035_ ( .A1(\EXU/CSRControl/_1162_ ), .A2(\EXU/CSRControl/_0253_ ), .ZN(\EXU/CSRControl/_1164_ ) );
AOI21_X1 \EXU/CSRControl/_2036_ ( .A(\EXU/CSRControl/_1374_ ), .B1(\EXU/CSRControl/_1163_ ), .B2(\EXU/CSRControl/_1164_ ), .ZN(\EXU/CSRControl/_0002_ ) );
INV_X1 \EXU/CSRControl/_2037_ ( .A(\EXU/CSRControl/_0304_ ), .ZN(\EXU/CSRControl/_1165_ ) );
BUF_X4 \EXU/CSRControl/_2038_ ( .A(\EXU/CSRControl/_1134_ ), .Z(\EXU/CSRControl/_1166_ ) );
NAND2_X1 \EXU/CSRControl/_2039_ ( .A1(\EXU/CSRControl/_1139_ ), .A2(\EXU/CSRControl/_0257_ ), .ZN(\EXU/CSRControl/_1167_ ) );
NAND3_X1 \EXU/CSRControl/_2040_ ( .A1(\EXU/CSRControl/_1150_ ), .A2(\EXU/CSRControl/_0193_ ), .A3(\EXU/CSRControl/_0809_ ), .ZN(\EXU/CSRControl/_1168_ ) );
NAND2_X1 \EXU/CSRControl/_2041_ ( .A1(\EXU/CSRControl/_1167_ ), .A2(\EXU/CSRControl/_1168_ ), .ZN(\EXU/CSRControl/_1169_ ) );
NAND3_X1 \EXU/CSRControl/_2042_ ( .A1(\EXU/CSRControl/_1143_ ), .A2(\EXU/CSRControl/_0826_ ), .A3(\EXU/CSRControl/_0161_ ), .ZN(\EXU/CSRControl/_1170_ ) );
NAND3_X1 \EXU/CSRControl/_2043_ ( .A1(\EXU/CSRControl/_1141_ ), .A2(\EXU/CSRControl/_0826_ ), .A3(\EXU/CSRControl/_0225_ ), .ZN(\EXU/CSRControl/_1171_ ) );
NAND2_X1 \EXU/CSRControl/_2044_ ( .A1(\EXU/CSRControl/_1170_ ), .A2(\EXU/CSRControl/_1171_ ), .ZN(\EXU/CSRControl/_1172_ ) );
OAI221_X1 \EXU/CSRControl/_2045_ ( .A(\EXU/CSRControl/_1135_ ), .B1(\EXU/CSRControl/_1165_ ), .B2(\EXU/CSRControl/_1166_ ), .C1(\EXU/CSRControl/_1169_ ), .C2(\EXU/CSRControl/_1172_ ), .ZN(\EXU/CSRControl/_1173_ ) );
CLKBUF_X2 \EXU/CSRControl/_2046_ ( .A(\EXU/CSRControl/_1154_ ), .Z(\EXU/CSRControl/_1174_ ) );
OR3_X1 \EXU/CSRControl/_2047_ ( .A1(\EXU/CSRControl/_1174_ ), .A2(\EXU/CSRControl/_0274_ ), .A3(\EXU/CSRControl/_1165_ ), .ZN(\EXU/CSRControl/_1175_ ) );
AND2_X1 \EXU/CSRControl/_2048_ ( .A1(\EXU/CSRControl/_1173_ ), .A2(\EXU/CSRControl/_1175_ ), .ZN(\EXU/CSRControl/_1176_ ) );
AOI21_X1 \EXU/CSRControl/_2049_ ( .A(\EXU/CSRControl/_0841_ ), .B1(\EXU/CSRControl/_1176_ ), .B2(\EXU/CSRControl/_1158_ ), .ZN(\EXU/CSRControl/_1177_ ) );
AOI211_X2 \EXU/CSRControl/_2050_ ( .A(\EXU/CSRControl/_1162_ ), .B(\EXU/CSRControl/_1177_ ), .C1(\EXU/CSRControl/_0253_ ), .C2(\EXU/CSRControl/_0841_ ), .ZN(\EXU/CSRControl/_1178_ ) );
NOR3_X1 \EXU/CSRControl/_2051_ ( .A1(\EXU/CSRControl/_1161_ ), .A2(\EXU/CSRControl/_0257_ ), .A3(\EXU/CSRControl/_0803_ ), .ZN(\EXU/CSRControl/_1179_ ) );
NOR3_X1 \EXU/CSRControl/_2052_ ( .A1(\EXU/CSRControl/_1178_ ), .A2(\EXU/CSRControl/_1374_ ), .A3(\EXU/CSRControl/_1179_ ), .ZN(\EXU/CSRControl/_0003_ ) );
AOI21_X1 \EXU/CSRControl/_2053_ ( .A(\EXU/CSRControl/_1374_ ), .B1(\EXU/CSRControl/_1162_ ), .B2(\EXU/CSRControl/_0230_ ), .ZN(\EXU/CSRControl/_1180_ ) );
BUF_X4 \EXU/CSRControl/_2054_ ( .A(\EXU/CSRControl/_1135_ ), .Z(\EXU/CSRControl/_1181_ ) );
INV_X1 \EXU/CSRControl/_2055_ ( .A(\EXU/CSRControl/_0277_ ), .ZN(\EXU/CSRControl/_1182_ ) );
BUF_X4 \EXU/CSRControl/_2056_ ( .A(\EXU/CSRControl/_1139_ ), .Z(\EXU/CSRControl/_1183_ ) );
NAND2_X1 \EXU/CSRControl/_2057_ ( .A1(\EXU/CSRControl/_1183_ ), .A2(\EXU/CSRControl/_0230_ ), .ZN(\EXU/CSRControl/_1184_ ) );
NAND2_X1 \EXU/CSRControl/_2058_ ( .A1(\EXU/CSRControl/_1149_ ), .A2(\EXU/CSRControl/_1184_ ), .ZN(\EXU/CSRControl/_1185_ ) );
BUF_X4 \EXU/CSRControl/_2059_ ( .A(\EXU/CSRControl/_1150_ ), .Z(\EXU/CSRControl/_1186_ ) );
BUF_X8 \EXU/CSRControl/_2060_ ( .A(\EXU/CSRControl/_1186_ ), .Z(\EXU/CSRControl/_1187_ ) );
BUF_X4 \EXU/CSRControl/_2061_ ( .A(\EXU/CSRControl/_0809_ ), .Z(\EXU/CSRControl/_1188_ ) );
BUF_X4 \EXU/CSRControl/_2062_ ( .A(\EXU/CSRControl/_1188_ ), .Z(\EXU/CSRControl/_1189_ ) );
NAND3_X1 \EXU/CSRControl/_2063_ ( .A1(\EXU/CSRControl/_1187_ ), .A2(\EXU/CSRControl/_0166_ ), .A3(\EXU/CSRControl/_1189_ ), .ZN(\EXU/CSRControl/_1190_ ) );
BUF_X4 \EXU/CSRControl/_2064_ ( .A(\EXU/CSRControl/_1141_ ), .Z(\EXU/CSRControl/_1191_ ) );
NAND3_X1 \EXU/CSRControl/_2065_ ( .A1(\EXU/CSRControl/_1191_ ), .A2(\EXU/CSRControl/_0827_ ), .A3(\EXU/CSRControl/_0198_ ), .ZN(\EXU/CSRControl/_1192_ ) );
BUF_X4 \EXU/CSRControl/_2066_ ( .A(\EXU/CSRControl/_1143_ ), .Z(\EXU/CSRControl/_1193_ ) );
NAND3_X1 \EXU/CSRControl/_2067_ ( .A1(\EXU/CSRControl/_1193_ ), .A2(\EXU/CSRControl/_0903_ ), .A3(\EXU/CSRControl/_0134_ ), .ZN(\EXU/CSRControl/_1194_ ) );
NAND3_X1 \EXU/CSRControl/_2068_ ( .A1(\EXU/CSRControl/_1190_ ), .A2(\EXU/CSRControl/_1192_ ), .A3(\EXU/CSRControl/_1194_ ), .ZN(\EXU/CSRControl/_1195_ ) );
OAI221_X1 \EXU/CSRControl/_2069_ ( .A(\EXU/CSRControl/_1181_ ), .B1(\EXU/CSRControl/_1182_ ), .B2(\EXU/CSRControl/_1166_ ), .C1(\EXU/CSRControl/_1185_ ), .C2(\EXU/CSRControl/_1195_ ), .ZN(\EXU/CSRControl/_1196_ ) );
OR3_X1 \EXU/CSRControl/_2070_ ( .A1(\EXU/CSRControl/_1174_ ), .A2(\EXU/CSRControl/_0274_ ), .A3(\EXU/CSRControl/_1182_ ), .ZN(\EXU/CSRControl/_1197_ ) );
AND2_X1 \EXU/CSRControl/_2071_ ( .A1(\EXU/CSRControl/_1196_ ), .A2(\EXU/CSRControl/_1197_ ), .ZN(\EXU/CSRControl/_1198_ ) );
NOR2_X1 \EXU/CSRControl/_2072_ ( .A1(\EXU/CSRControl/_1198_ ), .A2(\EXU/CSRControl/_1160_ ), .ZN(\EXU/CSRControl/_1199_ ) );
CLKBUF_X2 \EXU/CSRControl/_2073_ ( .A(\EXU/CSRControl/_0841_ ), .Z(\EXU/CSRControl/_1200_ ) );
AOI22_X1 \EXU/CSRControl/_2074_ ( .A1(\EXU/CSRControl/_1199_ ), .A2(\EXU/CSRControl/_1158_ ), .B1(\EXU/CSRControl/_1372_ ), .B2(\EXU/CSRControl/_1200_ ), .ZN(\EXU/CSRControl/_1201_ ) );
OAI21_X1 \EXU/CSRControl/_2075_ ( .A(\EXU/CSRControl/_1180_ ), .B1(\EXU/CSRControl/_1201_ ), .B2(\EXU/CSRControl/_1162_ ), .ZN(\EXU/CSRControl/_0004_ ) );
INV_X1 \EXU/CSRControl/_2076_ ( .A(\EXU/CSRControl/_1161_ ), .ZN(\EXU/CSRControl/_1202_ ) );
OR2_X2 \EXU/CSRControl/_2077_ ( .A1(\EXU/CSRControl/_1202_ ), .A2(\EXU/CSRControl/_0803_ ), .ZN(\EXU/CSRControl/_1203_ ) );
AND2_X4 \EXU/CSRControl/_2078_ ( .A1(\EXU/CSRControl/_1143_ ), .A2(\EXU/CSRControl/_0825_ ), .ZN(\EXU/CSRControl/_1204_ ) );
BUF_X4 \EXU/CSRControl/_2079_ ( .A(\EXU/CSRControl/_1204_ ), .Z(\EXU/CSRControl/_1205_ ) );
AOI22_X1 \EXU/CSRControl/_2080_ ( .A1(\EXU/CSRControl/_1205_ ), .A2(\EXU/CSRControl/_0135_ ), .B1(\EXU/CSRControl/_1183_ ), .B2(\EXU/CSRControl/_0231_ ), .ZN(\EXU/CSRControl/_1206_ ) );
BUF_X2 \EXU/CSRControl/_2081_ ( .A(\EXU/CSRControl/_1141_ ), .Z(\EXU/CSRControl/_1207_ ) );
BUF_X2 \EXU/CSRControl/_2082_ ( .A(\EXU/CSRControl/_0825_ ), .Z(\EXU/CSRControl/_1208_ ) );
AND3_X1 \EXU/CSRControl/_2083_ ( .A1(\EXU/CSRControl/_1207_ ), .A2(\EXU/CSRControl/_1208_ ), .A3(\EXU/CSRControl/_0199_ ), .ZN(\EXU/CSRControl/_1209_ ) );
NOR2_X1 \EXU/CSRControl/_2084_ ( .A1(\EXU/CSRControl/_1209_ ), .A2(\EXU/CSRControl/_1148_ ), .ZN(\EXU/CSRControl/_1210_ ) );
NAND3_X1 \EXU/CSRControl/_2085_ ( .A1(\EXU/CSRControl/_1187_ ), .A2(\EXU/CSRControl/_0167_ ), .A3(\EXU/CSRControl/_1189_ ), .ZN(\EXU/CSRControl/_1211_ ) );
NAND3_X1 \EXU/CSRControl/_2086_ ( .A1(\EXU/CSRControl/_1206_ ), .A2(\EXU/CSRControl/_1210_ ), .A3(\EXU/CSRControl/_1211_ ), .ZN(\EXU/CSRControl/_1212_ ) );
BUF_X4 \EXU/CSRControl/_2087_ ( .A(\EXU/CSRControl/_1135_ ), .Z(\EXU/CSRControl/_1213_ ) );
INV_X1 \EXU/CSRControl/_2088_ ( .A(\EXU/CSRControl/_0278_ ), .ZN(\EXU/CSRControl/_1214_ ) );
BUF_X4 \EXU/CSRControl/_2089_ ( .A(\EXU/CSRControl/_1166_ ), .Z(\EXU/CSRControl/_1215_ ) );
OAI211_X2 \EXU/CSRControl/_2090_ ( .A(\EXU/CSRControl/_1212_ ), .B(\EXU/CSRControl/_1213_ ), .C1(\EXU/CSRControl/_1214_ ), .C2(\EXU/CSRControl/_1215_ ), .ZN(\EXU/CSRControl/_1216_ ) );
OR3_X1 \EXU/CSRControl/_2091_ ( .A1(\EXU/CSRControl/_1174_ ), .A2(\EXU/CSRControl/_0274_ ), .A3(\EXU/CSRControl/_1214_ ), .ZN(\EXU/CSRControl/_1217_ ) );
AOI21_X1 \EXU/CSRControl/_2092_ ( .A(\EXU/CSRControl/_1203_ ), .B1(\EXU/CSRControl/_1216_ ), .B2(\EXU/CSRControl/_1217_ ), .ZN(\EXU/CSRControl/_1218_ ) );
AND2_X1 \EXU/CSRControl/_2093_ ( .A1(\EXU/CSRControl/_0841_ ), .A2(\EXU/CSRControl/_1373_ ), .ZN(\EXU/CSRControl/_1219_ ) );
MUX2_X1 \EXU/CSRControl/_2094_ ( .A(\EXU/CSRControl/_1219_ ), .B(\EXU/CSRControl/_0231_ ), .S(\EXU/CSRControl/_1162_ ), .Z(\EXU/CSRControl/_1220_ ) );
OR3_X1 \EXU/CSRControl/_2095_ ( .A1(\EXU/CSRControl/_1218_ ), .A2(\EXU/CSRControl/_1374_ ), .A3(\EXU/CSRControl/_1220_ ), .ZN(\EXU/CSRControl/_0005_ ) );
INV_X4 \EXU/CSRControl/_2096_ ( .A(\EXU/CSRControl/_1374_ ), .ZN(\EXU/CSRControl/_1221_ ) );
BUF_X4 \EXU/CSRControl/_2097_ ( .A(\EXU/CSRControl/_1221_ ), .Z(\EXU/CSRControl/_1222_ ) );
BUF_X4 \EXU/CSRControl/_2098_ ( .A(\EXU/CSRControl/_1222_ ), .Z(\EXU/CSRControl/_1223_ ) );
NAND3_X1 \EXU/CSRControl/_2099_ ( .A1(\EXU/CSRControl/_0803_ ), .A2(\EXU/CSRControl/_0272_ ), .A3(\EXU/CSRControl/_0230_ ), .ZN(\EXU/CSRControl/_1224_ ) );
OAI21_X1 \EXU/CSRControl/_2100_ ( .A(\EXU/CSRControl/_1372_ ), .B1(\EXU/CSRControl/_0801_ ), .B2(\EXU/CSRControl/_0273_ ), .ZN(\EXU/CSRControl/_1225_ ) );
NAND4_X1 \EXU/CSRControl/_2101_ ( .A1(\EXU/CSRControl/_0843_ ), .A2(\EXU/CSRControl/_1223_ ), .A3(\EXU/CSRControl/_1224_ ), .A4(\EXU/CSRControl/_1225_ ), .ZN(\EXU/CSRControl/_0006_ ) );
MUX2_X1 \EXU/CSRControl/_2102_ ( .A(\EXU/CSRControl/_1373_ ), .B(\EXU/CSRControl/_0231_ ), .S(\EXU/CSRControl/_0805_ ), .Z(\EXU/CSRControl/_1226_ ) );
OR3_X1 \EXU/CSRControl/_2103_ ( .A1(\EXU/CSRControl/_1226_ ), .A2(\EXU/CSRControl/_1374_ ), .A3(\EXU/CSRControl/_1200_ ), .ZN(\EXU/CSRControl/_0007_ ) );
NAND3_X1 \EXU/CSRControl/_2104_ ( .A1(\EXU/CSRControl/_0799_ ), .A2(\EXU/CSRControl/_0272_ ), .A3(\EXU/CSRControl/_0275_ ), .ZN(\EXU/CSRControl/_1227_ ) );
BUF_X4 \EXU/CSRControl/_2105_ ( .A(\EXU/CSRControl/_1143_ ), .Z(\EXU/CSRControl/_1228_ ) );
BUF_X4 \EXU/CSRControl/_2106_ ( .A(\EXU/CSRControl/_1208_ ), .Z(\EXU/CSRControl/_1229_ ) );
NAND3_X1 \EXU/CSRControl/_2107_ ( .A1(\EXU/CSRControl/_1228_ ), .A2(\EXU/CSRControl/_1229_ ), .A3(\EXU/CSRControl/_0132_ ), .ZN(\EXU/CSRControl/_1230_ ) );
BUF_X4 \EXU/CSRControl/_2108_ ( .A(\EXU/CSRControl/_1139_ ), .Z(\EXU/CSRControl/_1231_ ) );
NAND2_X1 \EXU/CSRControl/_2109_ ( .A1(\EXU/CSRControl/_1231_ ), .A2(\EXU/CSRControl/_0228_ ), .ZN(\EXU/CSRControl/_1232_ ) );
NAND2_X1 \EXU/CSRControl/_2110_ ( .A1(\EXU/CSRControl/_1230_ ), .A2(\EXU/CSRControl/_1232_ ), .ZN(\EXU/CSRControl/_1233_ ) );
BUF_X8 \EXU/CSRControl/_2111_ ( .A(\EXU/CSRControl/_1186_ ), .Z(\EXU/CSRControl/_1234_ ) );
BUF_X4 \EXU/CSRControl/_2112_ ( .A(\EXU/CSRControl/_1188_ ), .Z(\EXU/CSRControl/_1235_ ) );
NAND3_X1 \EXU/CSRControl/_2113_ ( .A1(\EXU/CSRControl/_1234_ ), .A2(\EXU/CSRControl/_0164_ ), .A3(\EXU/CSRControl/_1235_ ), .ZN(\EXU/CSRControl/_1236_ ) );
BUF_X4 \EXU/CSRControl/_2114_ ( .A(\EXU/CSRControl/_1207_ ), .Z(\EXU/CSRControl/_1237_ ) );
NAND3_X1 \EXU/CSRControl/_2115_ ( .A1(\EXU/CSRControl/_1237_ ), .A2(\EXU/CSRControl/_1229_ ), .A3(\EXU/CSRControl/_0196_ ), .ZN(\EXU/CSRControl/_1238_ ) );
NAND2_X1 \EXU/CSRControl/_2116_ ( .A1(\EXU/CSRControl/_1236_ ), .A2(\EXU/CSRControl/_1238_ ), .ZN(\EXU/CSRControl/_1239_ ) );
OAI211_X2 \EXU/CSRControl/_2117_ ( .A(\EXU/CSRControl/_1213_ ), .B(\EXU/CSRControl/_1227_ ), .C1(\EXU/CSRControl/_1233_ ), .C2(\EXU/CSRControl/_1239_ ), .ZN(\EXU/CSRControl/_1240_ ) );
NOR2_X2 \EXU/CSRControl/_2118_ ( .A1(\EXU/CSRControl/_1202_ ), .A2(\EXU/CSRControl/_0803_ ), .ZN(\EXU/CSRControl/_1241_ ) );
BUF_X2 \EXU/CSRControl/_2119_ ( .A(\EXU/CSRControl/_1241_ ), .Z(\EXU/CSRControl/_1242_ ) );
BUF_X8 \EXU/CSRControl/_2120_ ( .A(\EXU/CSRControl/_1242_ ), .Z(\EXU/CSRControl/_1243_ ) );
BUF_X4 \EXU/CSRControl/_2121_ ( .A(\EXU/CSRControl/_1155_ ), .Z(\EXU/CSRControl/_1244_ ) );
NAND2_X1 \EXU/CSRControl/_2122_ ( .A1(\EXU/CSRControl/_1244_ ), .A2(\EXU/CSRControl/_0275_ ), .ZN(\EXU/CSRControl/_1245_ ) );
AND3_X1 \EXU/CSRControl/_2123_ ( .A1(\EXU/CSRControl/_1240_ ), .A2(\EXU/CSRControl/_1243_ ), .A3(\EXU/CSRControl/_1245_ ), .ZN(\EXU/CSRControl/_1246_ ) );
BUF_X4 \EXU/CSRControl/_2124_ ( .A(\EXU/CSRControl/_1242_ ), .Z(\EXU/CSRControl/_1247_ ) );
OAI21_X1 \EXU/CSRControl/_2125_ ( .A(\EXU/CSRControl/_1223_ ), .B1(\EXU/CSRControl/_1247_ ), .B2(\EXU/CSRControl/_0228_ ), .ZN(\EXU/CSRControl/_1248_ ) );
NOR2_X1 \EXU/CSRControl/_2126_ ( .A1(\EXU/CSRControl/_1246_ ), .A2(\EXU/CSRControl/_1248_ ), .ZN(\EXU/CSRControl/_0008_ ) );
INV_X1 \EXU/CSRControl/_2127_ ( .A(\EXU/CSRControl/_0286_ ), .ZN(\EXU/CSRControl/_1249_ ) );
INV_X1 \EXU/CSRControl/_2128_ ( .A(\EXU/CSRControl/_0239_ ), .ZN(\EXU/CSRControl/_1250_ ) );
OR3_X1 \EXU/CSRControl/_2129_ ( .A1(\EXU/CSRControl/_1137_ ), .A2(\EXU/CSRControl/_1250_ ), .A3(\EXU/CSRControl/_1138_ ), .ZN(\EXU/CSRControl/_1251_ ) );
NAND3_X1 \EXU/CSRControl/_2130_ ( .A1(\EXU/CSRControl/_1186_ ), .A2(\EXU/CSRControl/_0175_ ), .A3(\EXU/CSRControl/_1188_ ), .ZN(\EXU/CSRControl/_1252_ ) );
NAND2_X1 \EXU/CSRControl/_2131_ ( .A1(\EXU/CSRControl/_1251_ ), .A2(\EXU/CSRControl/_1252_ ), .ZN(\EXU/CSRControl/_1253_ ) );
NAND3_X1 \EXU/CSRControl/_2132_ ( .A1(\EXU/CSRControl/_1193_ ), .A2(\EXU/CSRControl/_1117_ ), .A3(\EXU/CSRControl/_0143_ ), .ZN(\EXU/CSRControl/_1254_ ) );
NAND3_X1 \EXU/CSRControl/_2133_ ( .A1(\EXU/CSRControl/_1207_ ), .A2(\EXU/CSRControl/_1117_ ), .A3(\EXU/CSRControl/_0207_ ), .ZN(\EXU/CSRControl/_1255_ ) );
NAND2_X1 \EXU/CSRControl/_2134_ ( .A1(\EXU/CSRControl/_1254_ ), .A2(\EXU/CSRControl/_1255_ ), .ZN(\EXU/CSRControl/_1256_ ) );
OAI221_X1 \EXU/CSRControl/_2135_ ( .A(\EXU/CSRControl/_1181_ ), .B1(\EXU/CSRControl/_1249_ ), .B2(\EXU/CSRControl/_1166_ ), .C1(\EXU/CSRControl/_1253_ ), .C2(\EXU/CSRControl/_1256_ ), .ZN(\EXU/CSRControl/_1257_ ) );
OR3_X1 \EXU/CSRControl/_2136_ ( .A1(\EXU/CSRControl/_1174_ ), .A2(\EXU/CSRControl/_0274_ ), .A3(\EXU/CSRControl/_1249_ ), .ZN(\EXU/CSRControl/_1258_ ) );
AND3_X1 \EXU/CSRControl/_2137_ ( .A1(\EXU/CSRControl/_1257_ ), .A2(\EXU/CSRControl/_1242_ ), .A3(\EXU/CSRControl/_1258_ ), .ZN(\EXU/CSRControl/_1259_ ) );
AOI211_X2 \EXU/CSRControl/_2138_ ( .A(\EXU/CSRControl/_1374_ ), .B(\EXU/CSRControl/_1259_ ), .C1(\EXU/CSRControl/_1250_ ), .C2(\EXU/CSRControl/_1203_ ), .ZN(\EXU/CSRControl/_0009_ ) );
BUF_X4 \EXU/CSRControl/_2139_ ( .A(\EXU/CSRControl/_1221_ ), .Z(\EXU/CSRControl/_1260_ ) );
BUF_X4 \EXU/CSRControl/_2140_ ( .A(\EXU/CSRControl/_1242_ ), .Z(\EXU/CSRControl/_1261_ ) );
OAI21_X1 \EXU/CSRControl/_2141_ ( .A(\EXU/CSRControl/_1260_ ), .B1(\EXU/CSRControl/_1261_ ), .B2(\EXU/CSRControl/_0250_ ), .ZN(\EXU/CSRControl/_1262_ ) );
BUF_X4 \EXU/CSRControl/_2142_ ( .A(\EXU/CSRControl/_1135_ ), .Z(\EXU/CSRControl/_1263_ ) );
INV_X1 \EXU/CSRControl/_2143_ ( .A(\EXU/CSRControl/_0297_ ), .ZN(\EXU/CSRControl/_1264_ ) );
NAND2_X1 \EXU/CSRControl/_2144_ ( .A1(\EXU/CSRControl/_1231_ ), .A2(\EXU/CSRControl/_0250_ ), .ZN(\EXU/CSRControl/_1265_ ) );
NAND3_X1 \EXU/CSRControl/_2145_ ( .A1(\EXU/CSRControl/_1234_ ), .A2(\EXU/CSRControl/_0186_ ), .A3(\EXU/CSRControl/_1235_ ), .ZN(\EXU/CSRControl/_1266_ ) );
NAND2_X1 \EXU/CSRControl/_2146_ ( .A1(\EXU/CSRControl/_1265_ ), .A2(\EXU/CSRControl/_1266_ ), .ZN(\EXU/CSRControl/_1267_ ) );
NAND3_X1 \EXU/CSRControl/_2147_ ( .A1(\EXU/CSRControl/_1228_ ), .A2(\EXU/CSRControl/_1229_ ), .A3(\EXU/CSRControl/_0154_ ), .ZN(\EXU/CSRControl/_1268_ ) );
BUF_X4 \EXU/CSRControl/_2148_ ( .A(\EXU/CSRControl/_1208_ ), .Z(\EXU/CSRControl/_1269_ ) );
NAND3_X1 \EXU/CSRControl/_2149_ ( .A1(\EXU/CSRControl/_1237_ ), .A2(\EXU/CSRControl/_1269_ ), .A3(\EXU/CSRControl/_0218_ ), .ZN(\EXU/CSRControl/_1270_ ) );
NAND2_X1 \EXU/CSRControl/_2150_ ( .A1(\EXU/CSRControl/_1268_ ), .A2(\EXU/CSRControl/_1270_ ), .ZN(\EXU/CSRControl/_1271_ ) );
OAI221_X1 \EXU/CSRControl/_2151_ ( .A(\EXU/CSRControl/_1263_ ), .B1(\EXU/CSRControl/_1264_ ), .B2(\EXU/CSRControl/_1215_ ), .C1(\EXU/CSRControl/_1267_ ), .C2(\EXU/CSRControl/_1271_ ), .ZN(\EXU/CSRControl/_1272_ ) );
CLKBUF_X2 \EXU/CSRControl/_2152_ ( .A(\EXU/CSRControl/_1174_ ), .Z(\EXU/CSRControl/_1273_ ) );
OR3_X1 \EXU/CSRControl/_2153_ ( .A1(\EXU/CSRControl/_1273_ ), .A2(\EXU/CSRControl/_0274_ ), .A3(\EXU/CSRControl/_1264_ ), .ZN(\EXU/CSRControl/_1274_ ) );
AND2_X1 \EXU/CSRControl/_2154_ ( .A1(\EXU/CSRControl/_1272_ ), .A2(\EXU/CSRControl/_1274_ ), .ZN(\EXU/CSRControl/_1275_ ) );
BUF_X4 \EXU/CSRControl/_2155_ ( .A(\EXU/CSRControl/_1243_ ), .Z(\EXU/CSRControl/_1276_ ) );
AOI21_X1 \EXU/CSRControl/_2156_ ( .A(\EXU/CSRControl/_1262_ ), .B1(\EXU/CSRControl/_1275_ ), .B2(\EXU/CSRControl/_1276_ ), .ZN(\EXU/CSRControl/_0010_ ) );
OAI21_X1 \EXU/CSRControl/_2157_ ( .A(\EXU/CSRControl/_1260_ ), .B1(\EXU/CSRControl/_1261_ ), .B2(\EXU/CSRControl/_0254_ ), .ZN(\EXU/CSRControl/_1277_ ) );
AND2_X1 \EXU/CSRControl/_2158_ ( .A1(\EXU/CSRControl/_1141_ ), .A2(\EXU/CSRControl/_0825_ ), .ZN(\EXU/CSRControl/_1278_ ) );
AOI22_X1 \EXU/CSRControl/_2159_ ( .A1(\EXU/CSRControl/_1278_ ), .A2(\EXU/CSRControl/_0222_ ), .B1(\EXU/CSRControl/_1183_ ), .B2(\EXU/CSRControl/_0254_ ), .ZN(\EXU/CSRControl/_1279_ ) );
AND3_X1 \EXU/CSRControl/_2160_ ( .A1(\EXU/CSRControl/_1193_ ), .A2(\EXU/CSRControl/_0158_ ), .A3(\EXU/CSRControl/_1208_ ), .ZN(\EXU/CSRControl/_1280_ ) );
NOR2_X1 \EXU/CSRControl/_2161_ ( .A1(\EXU/CSRControl/_1280_ ), .A2(\EXU/CSRControl/_1148_ ), .ZN(\EXU/CSRControl/_1281_ ) );
NAND3_X1 \EXU/CSRControl/_2162_ ( .A1(\EXU/CSRControl/_1234_ ), .A2(\EXU/CSRControl/_0190_ ), .A3(\EXU/CSRControl/_1235_ ), .ZN(\EXU/CSRControl/_1282_ ) );
NAND3_X1 \EXU/CSRControl/_2163_ ( .A1(\EXU/CSRControl/_1279_ ), .A2(\EXU/CSRControl/_1281_ ), .A3(\EXU/CSRControl/_1282_ ), .ZN(\EXU/CSRControl/_1283_ ) );
NAND3_X1 \EXU/CSRControl/_2164_ ( .A1(\EXU/CSRControl/_0800_ ), .A2(\EXU/CSRControl/_0272_ ), .A3(\EXU/CSRControl/_0301_ ), .ZN(\EXU/CSRControl/_1284_ ) );
NAND3_X1 \EXU/CSRControl/_2165_ ( .A1(\EXU/CSRControl/_1283_ ), .A2(\EXU/CSRControl/_1213_ ), .A3(\EXU/CSRControl/_1284_ ), .ZN(\EXU/CSRControl/_1285_ ) );
NAND2_X1 \EXU/CSRControl/_2166_ ( .A1(\EXU/CSRControl/_1244_ ), .A2(\EXU/CSRControl/_0301_ ), .ZN(\EXU/CSRControl/_1286_ ) );
AND2_X1 \EXU/CSRControl/_2167_ ( .A1(\EXU/CSRControl/_1285_ ), .A2(\EXU/CSRControl/_1286_ ), .ZN(\EXU/CSRControl/_1287_ ) );
AOI21_X1 \EXU/CSRControl/_2168_ ( .A(\EXU/CSRControl/_1277_ ), .B1(\EXU/CSRControl/_1287_ ), .B2(\EXU/CSRControl/_1276_ ), .ZN(\EXU/CSRControl/_0011_ ) );
OAI21_X1 \EXU/CSRControl/_2169_ ( .A(\EXU/CSRControl/_1260_ ), .B1(\EXU/CSRControl/_1261_ ), .B2(\EXU/CSRControl/_0255_ ), .ZN(\EXU/CSRControl/_1288_ ) );
INV_X1 \EXU/CSRControl/_2170_ ( .A(\EXU/CSRControl/_0302_ ), .ZN(\EXU/CSRControl/_1289_ ) );
NAND2_X1 \EXU/CSRControl/_2171_ ( .A1(\EXU/CSRControl/_1231_ ), .A2(\EXU/CSRControl/_0255_ ), .ZN(\EXU/CSRControl/_1290_ ) );
NAND3_X1 \EXU/CSRControl/_2172_ ( .A1(\EXU/CSRControl/_1237_ ), .A2(\EXU/CSRControl/_1269_ ), .A3(\EXU/CSRControl/_0223_ ), .ZN(\EXU/CSRControl/_1291_ ) );
NAND3_X1 \EXU/CSRControl/_2173_ ( .A1(\EXU/CSRControl/_1228_ ), .A2(\EXU/CSRControl/_1269_ ), .A3(\EXU/CSRControl/_0159_ ), .ZN(\EXU/CSRControl/_1292_ ) );
NAND3_X1 \EXU/CSRControl/_2174_ ( .A1(\EXU/CSRControl/_1290_ ), .A2(\EXU/CSRControl/_1291_ ), .A3(\EXU/CSRControl/_1292_ ), .ZN(\EXU/CSRControl/_1293_ ) );
NAND3_X1 \EXU/CSRControl/_2175_ ( .A1(\EXU/CSRControl/_1187_ ), .A2(\EXU/CSRControl/_0191_ ), .A3(\EXU/CSRControl/_1189_ ), .ZN(\EXU/CSRControl/_1294_ ) );
NAND2_X1 \EXU/CSRControl/_2176_ ( .A1(\EXU/CSRControl/_1149_ ), .A2(\EXU/CSRControl/_1294_ ), .ZN(\EXU/CSRControl/_1295_ ) );
OAI221_X1 \EXU/CSRControl/_2177_ ( .A(\EXU/CSRControl/_1263_ ), .B1(\EXU/CSRControl/_1289_ ), .B2(\EXU/CSRControl/_1215_ ), .C1(\EXU/CSRControl/_1293_ ), .C2(\EXU/CSRControl/_1295_ ), .ZN(\EXU/CSRControl/_1296_ ) );
OR3_X1 \EXU/CSRControl/_2178_ ( .A1(\EXU/CSRControl/_1273_ ), .A2(\EXU/CSRControl/_0274_ ), .A3(\EXU/CSRControl/_1289_ ), .ZN(\EXU/CSRControl/_1297_ ) );
AND2_X1 \EXU/CSRControl/_2179_ ( .A1(\EXU/CSRControl/_1296_ ), .A2(\EXU/CSRControl/_1297_ ), .ZN(\EXU/CSRControl/_1298_ ) );
AOI21_X1 \EXU/CSRControl/_2180_ ( .A(\EXU/CSRControl/_1288_ ), .B1(\EXU/CSRControl/_1298_ ), .B2(\EXU/CSRControl/_1276_ ), .ZN(\EXU/CSRControl/_0012_ ) );
AND3_X1 \EXU/CSRControl/_2181_ ( .A1(\EXU/CSRControl/_1141_ ), .A2(\EXU/CSRControl/_0825_ ), .A3(\EXU/CSRControl/_0224_ ), .ZN(\EXU/CSRControl/_1299_ ) );
AOI21_X1 \EXU/CSRControl/_2182_ ( .A(\EXU/CSRControl/_1299_ ), .B1(\EXU/CSRControl/_0160_ ), .B2(\EXU/CSRControl/_1205_ ), .ZN(\EXU/CSRControl/_1300_ ) );
AND3_X1 \EXU/CSRControl/_2183_ ( .A1(\EXU/CSRControl/_1150_ ), .A2(\EXU/CSRControl/_0192_ ), .A3(\EXU/CSRControl/_0809_ ), .ZN(\EXU/CSRControl/_1301_ ) );
NOR2_X1 \EXU/CSRControl/_2184_ ( .A1(\EXU/CSRControl/_1301_ ), .A2(\EXU/CSRControl/_1148_ ), .ZN(\EXU/CSRControl/_1302_ ) );
INV_X1 \EXU/CSRControl/_2185_ ( .A(\EXU/CSRControl/_0256_ ), .ZN(\EXU/CSRControl/_1303_ ) );
OR3_X1 \EXU/CSRControl/_2186_ ( .A1(\EXU/CSRControl/_1137_ ), .A2(\EXU/CSRControl/_1303_ ), .A3(\EXU/CSRControl/_1138_ ), .ZN(\EXU/CSRControl/_1304_ ) );
NAND3_X1 \EXU/CSRControl/_2187_ ( .A1(\EXU/CSRControl/_1300_ ), .A2(\EXU/CSRControl/_1302_ ), .A3(\EXU/CSRControl/_1304_ ), .ZN(\EXU/CSRControl/_1305_ ) );
NAND3_X1 \EXU/CSRControl/_2188_ ( .A1(\EXU/CSRControl/_0799_ ), .A2(\EXU/CSRControl/_0272_ ), .A3(\EXU/CSRControl/_0303_ ), .ZN(\EXU/CSRControl/_1306_ ) );
NAND3_X1 \EXU/CSRControl/_2189_ ( .A1(\EXU/CSRControl/_1305_ ), .A2(\EXU/CSRControl/_1181_ ), .A3(\EXU/CSRControl/_1306_ ), .ZN(\EXU/CSRControl/_1307_ ) );
NAND2_X1 \EXU/CSRControl/_2190_ ( .A1(\EXU/CSRControl/_1244_ ), .A2(\EXU/CSRControl/_0303_ ), .ZN(\EXU/CSRControl/_1308_ ) );
AND3_X1 \EXU/CSRControl/_2191_ ( .A1(\EXU/CSRControl/_1307_ ), .A2(\EXU/CSRControl/_1242_ ), .A3(\EXU/CSRControl/_1308_ ), .ZN(\EXU/CSRControl/_1309_ ) );
AOI211_X2 \EXU/CSRControl/_2192_ ( .A(\EXU/CSRControl/_1374_ ), .B(\EXU/CSRControl/_1309_ ), .C1(\EXU/CSRControl/_1303_ ), .C2(\EXU/CSRControl/_1203_ ), .ZN(\EXU/CSRControl/_0013_ ) );
OAI21_X1 \EXU/CSRControl/_2193_ ( .A(\EXU/CSRControl/_1260_ ), .B1(\EXU/CSRControl/_1261_ ), .B2(\EXU/CSRControl/_0258_ ), .ZN(\EXU/CSRControl/_1310_ ) );
AND2_X4 \EXU/CSRControl/_2194_ ( .A1(\EXU/CSRControl/_1186_ ), .A2(\EXU/CSRControl/_1188_ ), .ZN(\EXU/CSRControl/_1311_ ) );
AOI22_X1 \EXU/CSRControl/_2195_ ( .A1(\EXU/CSRControl/_1311_ ), .A2(\EXU/CSRControl/_0194_ ), .B1(\EXU/CSRControl/_1205_ ), .B2(\EXU/CSRControl/_0162_ ), .ZN(\EXU/CSRControl/_1312_ ) );
AOI22_X1 \EXU/CSRControl/_2196_ ( .A1(\EXU/CSRControl/_1183_ ), .A2(\EXU/CSRControl/_0258_ ), .B1(\EXU/CSRControl/_1191_ ), .B2(\EXU/CSRControl/_1147_ ), .ZN(\EXU/CSRControl/_1313_ ) );
NAND3_X1 \EXU/CSRControl/_2197_ ( .A1(\EXU/CSRControl/_1237_ ), .A2(\EXU/CSRControl/_1229_ ), .A3(\EXU/CSRControl/_0226_ ), .ZN(\EXU/CSRControl/_1314_ ) );
NAND3_X1 \EXU/CSRControl/_2198_ ( .A1(\EXU/CSRControl/_1312_ ), .A2(\EXU/CSRControl/_1313_ ), .A3(\EXU/CSRControl/_1314_ ), .ZN(\EXU/CSRControl/_1315_ ) );
NAND3_X1 \EXU/CSRControl/_2199_ ( .A1(\EXU/CSRControl/_0799_ ), .A2(\EXU/CSRControl/_0272_ ), .A3(\EXU/CSRControl/_0305_ ), .ZN(\EXU/CSRControl/_1316_ ) );
NAND3_X1 \EXU/CSRControl/_2200_ ( .A1(\EXU/CSRControl/_1315_ ), .A2(\EXU/CSRControl/_1213_ ), .A3(\EXU/CSRControl/_1316_ ), .ZN(\EXU/CSRControl/_1317_ ) );
NAND2_X1 \EXU/CSRControl/_2201_ ( .A1(\EXU/CSRControl/_1244_ ), .A2(\EXU/CSRControl/_0305_ ), .ZN(\EXU/CSRControl/_1318_ ) );
AND2_X1 \EXU/CSRControl/_2202_ ( .A1(\EXU/CSRControl/_1317_ ), .A2(\EXU/CSRControl/_1318_ ), .ZN(\EXU/CSRControl/_1319_ ) );
AOI21_X1 \EXU/CSRControl/_2203_ ( .A(\EXU/CSRControl/_1310_ ), .B1(\EXU/CSRControl/_1319_ ), .B2(\EXU/CSRControl/_1276_ ), .ZN(\EXU/CSRControl/_0014_ ) );
NAND3_X1 \EXU/CSRControl/_2204_ ( .A1(\EXU/CSRControl/_0799_ ), .A2(\EXU/CSRControl/_0272_ ), .A3(\EXU/CSRControl/_0306_ ), .ZN(\EXU/CSRControl/_1320_ ) );
INV_X1 \EXU/CSRControl/_2205_ ( .A(\EXU/CSRControl/_0259_ ), .ZN(\EXU/CSRControl/_1321_ ) );
OR3_X1 \EXU/CSRControl/_2206_ ( .A1(\EXU/CSRControl/_1137_ ), .A2(\EXU/CSRControl/_1321_ ), .A3(\EXU/CSRControl/_1138_ ), .ZN(\EXU/CSRControl/_1322_ ) );
NAND3_X1 \EXU/CSRControl/_2207_ ( .A1(\EXU/CSRControl/_1186_ ), .A2(\EXU/CSRControl/_0195_ ), .A3(\EXU/CSRControl/_1188_ ), .ZN(\EXU/CSRControl/_1323_ ) );
NAND2_X1 \EXU/CSRControl/_2208_ ( .A1(\EXU/CSRControl/_1322_ ), .A2(\EXU/CSRControl/_1323_ ), .ZN(\EXU/CSRControl/_1324_ ) );
NAND3_X1 \EXU/CSRControl/_2209_ ( .A1(\EXU/CSRControl/_1193_ ), .A2(\EXU/CSRControl/_0874_ ), .A3(\EXU/CSRControl/_0163_ ), .ZN(\EXU/CSRControl/_1325_ ) );
NAND3_X1 \EXU/CSRControl/_2210_ ( .A1(\EXU/CSRControl/_1191_ ), .A2(\EXU/CSRControl/_1117_ ), .A3(\EXU/CSRControl/_0227_ ), .ZN(\EXU/CSRControl/_1326_ ) );
NAND2_X1 \EXU/CSRControl/_2211_ ( .A1(\EXU/CSRControl/_1325_ ), .A2(\EXU/CSRControl/_1326_ ), .ZN(\EXU/CSRControl/_1327_ ) );
OAI211_X2 \EXU/CSRControl/_2212_ ( .A(\EXU/CSRControl/_1181_ ), .B(\EXU/CSRControl/_1320_ ), .C1(\EXU/CSRControl/_1324_ ), .C2(\EXU/CSRControl/_1327_ ), .ZN(\EXU/CSRControl/_1328_ ) );
NAND2_X1 \EXU/CSRControl/_2213_ ( .A1(\EXU/CSRControl/_1244_ ), .A2(\EXU/CSRControl/_0306_ ), .ZN(\EXU/CSRControl/_1329_ ) );
AND3_X1 \EXU/CSRControl/_2214_ ( .A1(\EXU/CSRControl/_1328_ ), .A2(\EXU/CSRControl/_1242_ ), .A3(\EXU/CSRControl/_1329_ ), .ZN(\EXU/CSRControl/_1330_ ) );
AOI211_X2 \EXU/CSRControl/_2215_ ( .A(\EXU/CSRControl/_1374_ ), .B(\EXU/CSRControl/_1330_ ), .C1(\EXU/CSRControl/_1321_ ), .C2(\EXU/CSRControl/_1203_ ), .ZN(\EXU/CSRControl/_0015_ ) );
INV_X1 \EXU/CSRControl/_2216_ ( .A(\EXU/CSRControl/_0276_ ), .ZN(\EXU/CSRControl/_1331_ ) );
INV_X1 \EXU/CSRControl/_2217_ ( .A(\EXU/CSRControl/_0229_ ), .ZN(\EXU/CSRControl/_1332_ ) );
OR3_X1 \EXU/CSRControl/_2218_ ( .A1(\EXU/CSRControl/_1137_ ), .A2(\EXU/CSRControl/_1332_ ), .A3(\EXU/CSRControl/_1138_ ), .ZN(\EXU/CSRControl/_1333_ ) );
NAND3_X1 \EXU/CSRControl/_2219_ ( .A1(\EXU/CSRControl/_1186_ ), .A2(\EXU/CSRControl/_0165_ ), .A3(\EXU/CSRControl/_1188_ ), .ZN(\EXU/CSRControl/_1334_ ) );
NAND2_X1 \EXU/CSRControl/_2220_ ( .A1(\EXU/CSRControl/_1333_ ), .A2(\EXU/CSRControl/_1334_ ), .ZN(\EXU/CSRControl/_1335_ ) );
NAND3_X1 \EXU/CSRControl/_2221_ ( .A1(\EXU/CSRControl/_1193_ ), .A2(\EXU/CSRControl/_1117_ ), .A3(\EXU/CSRControl/_0133_ ), .ZN(\EXU/CSRControl/_1336_ ) );
NAND3_X1 \EXU/CSRControl/_2222_ ( .A1(\EXU/CSRControl/_1207_ ), .A2(\EXU/CSRControl/_1117_ ), .A3(\EXU/CSRControl/_0197_ ), .ZN(\EXU/CSRControl/_1337_ ) );
NAND2_X1 \EXU/CSRControl/_2223_ ( .A1(\EXU/CSRControl/_1336_ ), .A2(\EXU/CSRControl/_1337_ ), .ZN(\EXU/CSRControl/_1338_ ) );
OAI221_X1 \EXU/CSRControl/_2224_ ( .A(\EXU/CSRControl/_1181_ ), .B1(\EXU/CSRControl/_1331_ ), .B2(\EXU/CSRControl/_1166_ ), .C1(\EXU/CSRControl/_1335_ ), .C2(\EXU/CSRControl/_1338_ ), .ZN(\EXU/CSRControl/_1339_ ) );
OR3_X1 \EXU/CSRControl/_2225_ ( .A1(\EXU/CSRControl/_1174_ ), .A2(\EXU/CSRControl/_0274_ ), .A3(\EXU/CSRControl/_1331_ ), .ZN(\EXU/CSRControl/_1340_ ) );
AND3_X1 \EXU/CSRControl/_2226_ ( .A1(\EXU/CSRControl/_1339_ ), .A2(\EXU/CSRControl/_1242_ ), .A3(\EXU/CSRControl/_1340_ ), .ZN(\EXU/CSRControl/_1341_ ) );
AOI211_X2 \EXU/CSRControl/_2227_ ( .A(\EXU/CSRControl/_1374_ ), .B(\EXU/CSRControl/_1341_ ), .C1(\EXU/CSRControl/_1332_ ), .C2(\EXU/CSRControl/_1203_ ), .ZN(\EXU/CSRControl/_0016_ ) );
INV_X1 \EXU/CSRControl/_2228_ ( .A(\EXU/CSRControl/_0279_ ), .ZN(\EXU/CSRControl/_1342_ ) );
NAND2_X1 \EXU/CSRControl/_2229_ ( .A1(\EXU/CSRControl/_1231_ ), .A2(\EXU/CSRControl/_0232_ ), .ZN(\EXU/CSRControl/_1343_ ) );
NAND2_X1 \EXU/CSRControl/_2230_ ( .A1(\EXU/CSRControl/_1149_ ), .A2(\EXU/CSRControl/_1343_ ), .ZN(\EXU/CSRControl/_1344_ ) );
NAND3_X1 \EXU/CSRControl/_2231_ ( .A1(\EXU/CSRControl/_1187_ ), .A2(\EXU/CSRControl/_0168_ ), .A3(\EXU/CSRControl/_1189_ ), .ZN(\EXU/CSRControl/_1345_ ) );
NAND3_X1 \EXU/CSRControl/_2232_ ( .A1(\EXU/CSRControl/_1191_ ), .A2(\EXU/CSRControl/_0827_ ), .A3(\EXU/CSRControl/_0200_ ), .ZN(\EXU/CSRControl/_1346_ ) );
NAND3_X1 \EXU/CSRControl/_2233_ ( .A1(\EXU/CSRControl/_1193_ ), .A2(\EXU/CSRControl/_0827_ ), .A3(\EXU/CSRControl/_0136_ ), .ZN(\EXU/CSRControl/_1347_ ) );
NAND3_X1 \EXU/CSRControl/_2234_ ( .A1(\EXU/CSRControl/_1345_ ), .A2(\EXU/CSRControl/_1346_ ), .A3(\EXU/CSRControl/_1347_ ), .ZN(\EXU/CSRControl/_1348_ ) );
OAI221_X1 \EXU/CSRControl/_2235_ ( .A(\EXU/CSRControl/_1263_ ), .B1(\EXU/CSRControl/_1342_ ), .B2(\EXU/CSRControl/_1215_ ), .C1(\EXU/CSRControl/_1344_ ), .C2(\EXU/CSRControl/_1348_ ), .ZN(\EXU/CSRControl/_1349_ ) );
OR3_X1 \EXU/CSRControl/_2236_ ( .A1(\EXU/CSRControl/_1273_ ), .A2(\EXU/CSRControl/_0274_ ), .A3(\EXU/CSRControl/_1342_ ), .ZN(\EXU/CSRControl/_1350_ ) );
AND3_X1 \EXU/CSRControl/_2237_ ( .A1(\EXU/CSRControl/_1349_ ), .A2(\EXU/CSRControl/_1243_ ), .A3(\EXU/CSRControl/_1350_ ), .ZN(\EXU/CSRControl/_1351_ ) );
OAI21_X1 \EXU/CSRControl/_2238_ ( .A(\EXU/CSRControl/_1223_ ), .B1(\EXU/CSRControl/_1247_ ), .B2(\EXU/CSRControl/_0232_ ), .ZN(\EXU/CSRControl/_1352_ ) );
NOR2_X1 \EXU/CSRControl/_2239_ ( .A1(\EXU/CSRControl/_1351_ ), .A2(\EXU/CSRControl/_1352_ ), .ZN(\EXU/CSRControl/_0017_ ) );
OAI21_X1 \EXU/CSRControl/_2240_ ( .A(\EXU/CSRControl/_1260_ ), .B1(\EXU/CSRControl/_1261_ ), .B2(\EXU/CSRControl/_0233_ ), .ZN(\EXU/CSRControl/_1353_ ) );
AOI22_X1 \EXU/CSRControl/_2241_ ( .A1(\EXU/CSRControl/_1311_ ), .A2(\EXU/CSRControl/_0169_ ), .B1(\EXU/CSRControl/_1205_ ), .B2(\EXU/CSRControl/_0137_ ), .ZN(\EXU/CSRControl/_1354_ ) );
AOI22_X1 \EXU/CSRControl/_2242_ ( .A1(\EXU/CSRControl/_1183_ ), .A2(\EXU/CSRControl/_0233_ ), .B1(\EXU/CSRControl/_1191_ ), .B2(\EXU/CSRControl/_1147_ ), .ZN(\EXU/CSRControl/_1355_ ) );
NAND3_X1 \EXU/CSRControl/_2243_ ( .A1(\EXU/CSRControl/_1237_ ), .A2(\EXU/CSRControl/_1229_ ), .A3(\EXU/CSRControl/_0201_ ), .ZN(\EXU/CSRControl/_1356_ ) );
NAND3_X1 \EXU/CSRControl/_2244_ ( .A1(\EXU/CSRControl/_1354_ ), .A2(\EXU/CSRControl/_1355_ ), .A3(\EXU/CSRControl/_1356_ ), .ZN(\EXU/CSRControl/_1357_ ) );
NAND3_X1 \EXU/CSRControl/_2245_ ( .A1(\EXU/CSRControl/_0799_ ), .A2(\EXU/CSRControl/_0272_ ), .A3(\EXU/CSRControl/_0280_ ), .ZN(\EXU/CSRControl/_1358_ ) );
NAND3_X1 \EXU/CSRControl/_2246_ ( .A1(\EXU/CSRControl/_1357_ ), .A2(\EXU/CSRControl/_1213_ ), .A3(\EXU/CSRControl/_1358_ ), .ZN(\EXU/CSRControl/_1359_ ) );
NAND2_X1 \EXU/CSRControl/_2247_ ( .A1(\EXU/CSRControl/_1244_ ), .A2(\EXU/CSRControl/_0280_ ), .ZN(\EXU/CSRControl/_1360_ ) );
AND2_X1 \EXU/CSRControl/_2248_ ( .A1(\EXU/CSRControl/_1359_ ), .A2(\EXU/CSRControl/_1360_ ), .ZN(\EXU/CSRControl/_1361_ ) );
AOI21_X1 \EXU/CSRControl/_2249_ ( .A(\EXU/CSRControl/_1353_ ), .B1(\EXU/CSRControl/_1361_ ), .B2(\EXU/CSRControl/_1276_ ), .ZN(\EXU/CSRControl/_0018_ ) );
INV_X1 \EXU/CSRControl/_2250_ ( .A(\EXU/CSRControl/_0281_ ), .ZN(\EXU/CSRControl/_1362_ ) );
NAND2_X1 \EXU/CSRControl/_2251_ ( .A1(\EXU/CSRControl/_1231_ ), .A2(\EXU/CSRControl/_0234_ ), .ZN(\EXU/CSRControl/_1363_ ) );
NAND3_X1 \EXU/CSRControl/_2252_ ( .A1(\EXU/CSRControl/_1234_ ), .A2(\EXU/CSRControl/_0170_ ), .A3(\EXU/CSRControl/_1235_ ), .ZN(\EXU/CSRControl/_1364_ ) );
NAND2_X1 \EXU/CSRControl/_2253_ ( .A1(\EXU/CSRControl/_1363_ ), .A2(\EXU/CSRControl/_1364_ ), .ZN(\EXU/CSRControl/_1365_ ) );
NAND3_X1 \EXU/CSRControl/_2254_ ( .A1(\EXU/CSRControl/_1228_ ), .A2(\EXU/CSRControl/_1229_ ), .A3(\EXU/CSRControl/_0138_ ), .ZN(\EXU/CSRControl/_1366_ ) );
NAND3_X1 \EXU/CSRControl/_2255_ ( .A1(\EXU/CSRControl/_1237_ ), .A2(\EXU/CSRControl/_1269_ ), .A3(\EXU/CSRControl/_0202_ ), .ZN(\EXU/CSRControl/_1367_ ) );
NAND2_X1 \EXU/CSRControl/_2256_ ( .A1(\EXU/CSRControl/_1366_ ), .A2(\EXU/CSRControl/_1367_ ), .ZN(\EXU/CSRControl/_1368_ ) );
OAI221_X1 \EXU/CSRControl/_2257_ ( .A(\EXU/CSRControl/_1263_ ), .B1(\EXU/CSRControl/_1362_ ), .B2(\EXU/CSRControl/_1215_ ), .C1(\EXU/CSRControl/_1365_ ), .C2(\EXU/CSRControl/_1368_ ), .ZN(\EXU/CSRControl/_1369_ ) );
OR3_X1 \EXU/CSRControl/_2258_ ( .A1(\EXU/CSRControl/_1273_ ), .A2(\EXU/CSRControl/_0274_ ), .A3(\EXU/CSRControl/_1362_ ), .ZN(\EXU/CSRControl/_1370_ ) );
AND3_X1 \EXU/CSRControl/_2259_ ( .A1(\EXU/CSRControl/_1369_ ), .A2(\EXU/CSRControl/_1243_ ), .A3(\EXU/CSRControl/_1370_ ), .ZN(\EXU/CSRControl/_1371_ ) );
OAI21_X1 \EXU/CSRControl/_2260_ ( .A(\EXU/CSRControl/_1223_ ), .B1(\EXU/CSRControl/_1247_ ), .B2(\EXU/CSRControl/_0234_ ), .ZN(\EXU/CSRControl/_0371_ ) );
NOR2_X1 \EXU/CSRControl/_2261_ ( .A1(\EXU/CSRControl/_1371_ ), .A2(\EXU/CSRControl/_0371_ ), .ZN(\EXU/CSRControl/_0019_ ) );
OAI21_X1 \EXU/CSRControl/_2262_ ( .A(\EXU/CSRControl/_1260_ ), .B1(\EXU/CSRControl/_1261_ ), .B2(\EXU/CSRControl/_0235_ ), .ZN(\EXU/CSRControl/_0372_ ) );
INV_X1 \EXU/CSRControl/_2263_ ( .A(\EXU/CSRControl/_0282_ ), .ZN(\EXU/CSRControl/_0373_ ) );
NAND2_X1 \EXU/CSRControl/_2264_ ( .A1(\EXU/CSRControl/_1231_ ), .A2(\EXU/CSRControl/_0235_ ), .ZN(\EXU/CSRControl/_0374_ ) );
NAND3_X1 \EXU/CSRControl/_2265_ ( .A1(\EXU/CSRControl/_1237_ ), .A2(\EXU/CSRControl/_1269_ ), .A3(\EXU/CSRControl/_0203_ ), .ZN(\EXU/CSRControl/_0375_ ) );
NAND3_X1 \EXU/CSRControl/_2266_ ( .A1(\EXU/CSRControl/_1228_ ), .A2(\EXU/CSRControl/_0827_ ), .A3(\EXU/CSRControl/_0139_ ), .ZN(\EXU/CSRControl/_0376_ ) );
NAND3_X1 \EXU/CSRControl/_2267_ ( .A1(\EXU/CSRControl/_0374_ ), .A2(\EXU/CSRControl/_0375_ ), .A3(\EXU/CSRControl/_0376_ ), .ZN(\EXU/CSRControl/_0377_ ) );
NAND3_X1 \EXU/CSRControl/_2268_ ( .A1(\EXU/CSRControl/_1187_ ), .A2(\EXU/CSRControl/_0171_ ), .A3(\EXU/CSRControl/_1189_ ), .ZN(\EXU/CSRControl/_0378_ ) );
NAND2_X1 \EXU/CSRControl/_2269_ ( .A1(\EXU/CSRControl/_1149_ ), .A2(\EXU/CSRControl/_0378_ ), .ZN(\EXU/CSRControl/_0379_ ) );
OAI221_X1 \EXU/CSRControl/_2270_ ( .A(\EXU/CSRControl/_1263_ ), .B1(\EXU/CSRControl/_0373_ ), .B2(\EXU/CSRControl/_1166_ ), .C1(\EXU/CSRControl/_0377_ ), .C2(\EXU/CSRControl/_0379_ ), .ZN(\EXU/CSRControl/_0380_ ) );
OR3_X1 \EXU/CSRControl/_2271_ ( .A1(\EXU/CSRControl/_1273_ ), .A2(\EXU/CSRControl/_0274_ ), .A3(\EXU/CSRControl/_0373_ ), .ZN(\EXU/CSRControl/_0381_ ) );
AND2_X1 \EXU/CSRControl/_2272_ ( .A1(\EXU/CSRControl/_0380_ ), .A2(\EXU/CSRControl/_0381_ ), .ZN(\EXU/CSRControl/_0382_ ) );
AOI21_X1 \EXU/CSRControl/_2273_ ( .A(\EXU/CSRControl/_0372_ ), .B1(\EXU/CSRControl/_0382_ ), .B2(\EXU/CSRControl/_1276_ ), .ZN(\EXU/CSRControl/_0020_ ) );
NAND3_X1 \EXU/CSRControl/_2274_ ( .A1(\EXU/CSRControl/_0799_ ), .A2(\EXU/CSRControl/_0272_ ), .A3(\EXU/CSRControl/_0283_ ), .ZN(\EXU/CSRControl/_0383_ ) );
INV_X1 \EXU/CSRControl/_2275_ ( .A(\EXU/CSRControl/_0236_ ), .ZN(\EXU/CSRControl/_0384_ ) );
OR3_X1 \EXU/CSRControl/_2276_ ( .A1(\EXU/CSRControl/_1137_ ), .A2(\EXU/CSRControl/_0384_ ), .A3(\EXU/CSRControl/_1138_ ), .ZN(\EXU/CSRControl/_0385_ ) );
NAND3_X1 \EXU/CSRControl/_2277_ ( .A1(\EXU/CSRControl/_1193_ ), .A2(\EXU/CSRControl/_1117_ ), .A3(\EXU/CSRControl/_0140_ ), .ZN(\EXU/CSRControl/_0386_ ) );
NAND3_X1 \EXU/CSRControl/_2278_ ( .A1(\EXU/CSRControl/_1186_ ), .A2(\EXU/CSRControl/_0172_ ), .A3(\EXU/CSRControl/_1188_ ), .ZN(\EXU/CSRControl/_0387_ ) );
NAND3_X1 \EXU/CSRControl/_2279_ ( .A1(\EXU/CSRControl/_0385_ ), .A2(\EXU/CSRControl/_0386_ ), .A3(\EXU/CSRControl/_0387_ ), .ZN(\EXU/CSRControl/_0388_ ) );
NAND3_X1 \EXU/CSRControl/_2280_ ( .A1(\EXU/CSRControl/_1191_ ), .A2(\EXU/CSRControl/_1117_ ), .A3(\EXU/CSRControl/_0204_ ), .ZN(\EXU/CSRControl/_0389_ ) );
NAND2_X1 \EXU/CSRControl/_2281_ ( .A1(\EXU/CSRControl/_1149_ ), .A2(\EXU/CSRControl/_0389_ ), .ZN(\EXU/CSRControl/_0390_ ) );
OAI211_X2 \EXU/CSRControl/_2282_ ( .A(\EXU/CSRControl/_1181_ ), .B(\EXU/CSRControl/_0383_ ), .C1(\EXU/CSRControl/_0388_ ), .C2(\EXU/CSRControl/_0390_ ), .ZN(\EXU/CSRControl/_0391_ ) );
NAND2_X1 \EXU/CSRControl/_2283_ ( .A1(\EXU/CSRControl/_1155_ ), .A2(\EXU/CSRControl/_0283_ ), .ZN(\EXU/CSRControl/_0392_ ) );
AND3_X1 \EXU/CSRControl/_2284_ ( .A1(\EXU/CSRControl/_0391_ ), .A2(\EXU/CSRControl/_1242_ ), .A3(\EXU/CSRControl/_0392_ ), .ZN(\EXU/CSRControl/_0393_ ) );
AOI211_X2 \EXU/CSRControl/_2285_ ( .A(\EXU/CSRControl/_1374_ ), .B(\EXU/CSRControl/_0393_ ), .C1(\EXU/CSRControl/_0384_ ), .C2(\EXU/CSRControl/_1203_ ), .ZN(\EXU/CSRControl/_0021_ ) );
INV_X1 \EXU/CSRControl/_2286_ ( .A(\EXU/CSRControl/_0284_ ), .ZN(\EXU/CSRControl/_0394_ ) );
INV_X1 \EXU/CSRControl/_2287_ ( .A(\EXU/CSRControl/_0237_ ), .ZN(\EXU/CSRControl/_0395_ ) );
OR3_X1 \EXU/CSRControl/_2288_ ( .A1(\EXU/CSRControl/_1137_ ), .A2(\EXU/CSRControl/_0395_ ), .A3(\EXU/CSRControl/_1138_ ), .ZN(\EXU/CSRControl/_0396_ ) );
NAND3_X1 \EXU/CSRControl/_2289_ ( .A1(\EXU/CSRControl/_1186_ ), .A2(\EXU/CSRControl/_0173_ ), .A3(\EXU/CSRControl/_1188_ ), .ZN(\EXU/CSRControl/_0397_ ) );
NAND2_X1 \EXU/CSRControl/_2290_ ( .A1(\EXU/CSRControl/_0396_ ), .A2(\EXU/CSRControl/_0397_ ), .ZN(\EXU/CSRControl/_0398_ ) );
NAND3_X1 \EXU/CSRControl/_2291_ ( .A1(\EXU/CSRControl/_1193_ ), .A2(\EXU/CSRControl/_1117_ ), .A3(\EXU/CSRControl/_0141_ ), .ZN(\EXU/CSRControl/_0399_ ) );
NAND3_X1 \EXU/CSRControl/_2292_ ( .A1(\EXU/CSRControl/_1207_ ), .A2(\EXU/CSRControl/_1208_ ), .A3(\EXU/CSRControl/_0205_ ), .ZN(\EXU/CSRControl/_0400_ ) );
NAND2_X1 \EXU/CSRControl/_2293_ ( .A1(\EXU/CSRControl/_0399_ ), .A2(\EXU/CSRControl/_0400_ ), .ZN(\EXU/CSRControl/_0401_ ) );
OAI221_X1 \EXU/CSRControl/_2294_ ( .A(\EXU/CSRControl/_1181_ ), .B1(\EXU/CSRControl/_0394_ ), .B2(\EXU/CSRControl/_1166_ ), .C1(\EXU/CSRControl/_0398_ ), .C2(\EXU/CSRControl/_0401_ ), .ZN(\EXU/CSRControl/_0402_ ) );
OR3_X1 \EXU/CSRControl/_2295_ ( .A1(\EXU/CSRControl/_1174_ ), .A2(\EXU/CSRControl/_0274_ ), .A3(\EXU/CSRControl/_0394_ ), .ZN(\EXU/CSRControl/_0403_ ) );
AND3_X1 \EXU/CSRControl/_2296_ ( .A1(\EXU/CSRControl/_0402_ ), .A2(\EXU/CSRControl/_1242_ ), .A3(\EXU/CSRControl/_0403_ ), .ZN(\EXU/CSRControl/_0404_ ) );
AOI211_X2 \EXU/CSRControl/_2297_ ( .A(\EXU/CSRControl/_1374_ ), .B(\EXU/CSRControl/_0404_ ), .C1(\EXU/CSRControl/_0395_ ), .C2(\EXU/CSRControl/_1203_ ), .ZN(\EXU/CSRControl/_0022_ ) );
OAI21_X1 \EXU/CSRControl/_2298_ ( .A(\EXU/CSRControl/_1260_ ), .B1(\EXU/CSRControl/_1261_ ), .B2(\EXU/CSRControl/_0238_ ), .ZN(\EXU/CSRControl/_0405_ ) );
INV_X1 \EXU/CSRControl/_2299_ ( .A(\EXU/CSRControl/_0285_ ), .ZN(\EXU/CSRControl/_0406_ ) );
NAND2_X1 \EXU/CSRControl/_2300_ ( .A1(\EXU/CSRControl/_1231_ ), .A2(\EXU/CSRControl/_0238_ ), .ZN(\EXU/CSRControl/_0407_ ) );
NAND3_X1 \EXU/CSRControl/_2301_ ( .A1(\EXU/CSRControl/_1228_ ), .A2(\EXU/CSRControl/_1229_ ), .A3(\EXU/CSRControl/_0142_ ), .ZN(\EXU/CSRControl/_0408_ ) );
NAND2_X1 \EXU/CSRControl/_2302_ ( .A1(\EXU/CSRControl/_0407_ ), .A2(\EXU/CSRControl/_0408_ ), .ZN(\EXU/CSRControl/_0409_ ) );
NAND3_X2 \EXU/CSRControl/_2303_ ( .A1(\EXU/CSRControl/_1234_ ), .A2(\EXU/CSRControl/_0174_ ), .A3(\EXU/CSRControl/_1235_ ), .ZN(\EXU/CSRControl/_0410_ ) );
NAND3_X1 \EXU/CSRControl/_2304_ ( .A1(\EXU/CSRControl/_1191_ ), .A2(\EXU/CSRControl/_1269_ ), .A3(\EXU/CSRControl/_0206_ ), .ZN(\EXU/CSRControl/_0411_ ) );
NAND2_X1 \EXU/CSRControl/_2305_ ( .A1(\EXU/CSRControl/_0410_ ), .A2(\EXU/CSRControl/_0411_ ), .ZN(\EXU/CSRControl/_0412_ ) );
OAI221_X1 \EXU/CSRControl/_2306_ ( .A(\EXU/CSRControl/_1263_ ), .B1(\EXU/CSRControl/_0406_ ), .B2(\EXU/CSRControl/_1166_ ), .C1(\EXU/CSRControl/_0409_ ), .C2(\EXU/CSRControl/_0412_ ), .ZN(\EXU/CSRControl/_0413_ ) );
OR3_X1 \EXU/CSRControl/_2307_ ( .A1(\EXU/CSRControl/_1273_ ), .A2(\EXU/CSRControl/_0274_ ), .A3(\EXU/CSRControl/_0406_ ), .ZN(\EXU/CSRControl/_0414_ ) );
AND2_X1 \EXU/CSRControl/_2308_ ( .A1(\EXU/CSRControl/_0413_ ), .A2(\EXU/CSRControl/_0414_ ), .ZN(\EXU/CSRControl/_0415_ ) );
AOI21_X1 \EXU/CSRControl/_2309_ ( .A(\EXU/CSRControl/_0405_ ), .B1(\EXU/CSRControl/_0415_ ), .B2(\EXU/CSRControl/_1276_ ), .ZN(\EXU/CSRControl/_0023_ ) );
OAI21_X1 \EXU/CSRControl/_2310_ ( .A(\EXU/CSRControl/_1260_ ), .B1(\EXU/CSRControl/_1261_ ), .B2(\EXU/CSRControl/_0240_ ), .ZN(\EXU/CSRControl/_0416_ ) );
INV_X1 \EXU/CSRControl/_2311_ ( .A(\EXU/CSRControl/_0287_ ), .ZN(\EXU/CSRControl/_0417_ ) );
NAND2_X1 \EXU/CSRControl/_2312_ ( .A1(\EXU/CSRControl/_1183_ ), .A2(\EXU/CSRControl/_0240_ ), .ZN(\EXU/CSRControl/_0418_ ) );
NAND3_X1 \EXU/CSRControl/_2313_ ( .A1(\EXU/CSRControl/_1187_ ), .A2(\EXU/CSRControl/_0176_ ), .A3(\EXU/CSRControl/_1189_ ), .ZN(\EXU/CSRControl/_0419_ ) );
NAND3_X1 \EXU/CSRControl/_2314_ ( .A1(\EXU/CSRControl/_1191_ ), .A2(\EXU/CSRControl/_0827_ ), .A3(\EXU/CSRControl/_0208_ ), .ZN(\EXU/CSRControl/_0420_ ) );
NAND3_X1 \EXU/CSRControl/_2315_ ( .A1(\EXU/CSRControl/_0418_ ), .A2(\EXU/CSRControl/_0419_ ), .A3(\EXU/CSRControl/_0420_ ), .ZN(\EXU/CSRControl/_0421_ ) );
NAND3_X1 \EXU/CSRControl/_2316_ ( .A1(\EXU/CSRControl/_1228_ ), .A2(\EXU/CSRControl/_1269_ ), .A3(\EXU/CSRControl/_0144_ ), .ZN(\EXU/CSRControl/_0422_ ) );
NAND2_X1 \EXU/CSRControl/_2317_ ( .A1(\EXU/CSRControl/_1149_ ), .A2(\EXU/CSRControl/_0422_ ), .ZN(\EXU/CSRControl/_0423_ ) );
OAI221_X1 \EXU/CSRControl/_2318_ ( .A(\EXU/CSRControl/_1181_ ), .B1(\EXU/CSRControl/_0417_ ), .B2(\EXU/CSRControl/_1166_ ), .C1(\EXU/CSRControl/_0421_ ), .C2(\EXU/CSRControl/_0423_ ), .ZN(\EXU/CSRControl/_0424_ ) );
OR3_X1 \EXU/CSRControl/_2319_ ( .A1(\EXU/CSRControl/_1273_ ), .A2(\EXU/CSRControl/_0274_ ), .A3(\EXU/CSRControl/_0417_ ), .ZN(\EXU/CSRControl/_0425_ ) );
AND2_X1 \EXU/CSRControl/_2320_ ( .A1(\EXU/CSRControl/_0424_ ), .A2(\EXU/CSRControl/_0425_ ), .ZN(\EXU/CSRControl/_0426_ ) );
AOI21_X1 \EXU/CSRControl/_2321_ ( .A(\EXU/CSRControl/_0416_ ), .B1(\EXU/CSRControl/_0426_ ), .B2(\EXU/CSRControl/_1276_ ), .ZN(\EXU/CSRControl/_0024_ ) );
OAI21_X1 \EXU/CSRControl/_2322_ ( .A(\EXU/CSRControl/_1260_ ), .B1(\EXU/CSRControl/_1261_ ), .B2(\EXU/CSRControl/_0241_ ), .ZN(\EXU/CSRControl/_0427_ ) );
AOI22_X1 \EXU/CSRControl/_2323_ ( .A1(\EXU/CSRControl/_1278_ ), .A2(\EXU/CSRControl/_0209_ ), .B1(\EXU/CSRControl/_1183_ ), .B2(\EXU/CSRControl/_0241_ ), .ZN(\EXU/CSRControl/_0428_ ) );
AND3_X1 \EXU/CSRControl/_2324_ ( .A1(\EXU/CSRControl/_1143_ ), .A2(\EXU/CSRControl/_0145_ ), .A3(\EXU/CSRControl/_0826_ ), .ZN(\EXU/CSRControl/_0429_ ) );
NOR2_X1 \EXU/CSRControl/_2325_ ( .A1(\EXU/CSRControl/_0429_ ), .A2(\EXU/CSRControl/_1148_ ), .ZN(\EXU/CSRControl/_0430_ ) );
NAND3_X1 \EXU/CSRControl/_2326_ ( .A1(\EXU/CSRControl/_1187_ ), .A2(\EXU/CSRControl/_0177_ ), .A3(\EXU/CSRControl/_1189_ ), .ZN(\EXU/CSRControl/_0431_ ) );
NAND3_X1 \EXU/CSRControl/_2327_ ( .A1(\EXU/CSRControl/_0428_ ), .A2(\EXU/CSRControl/_0430_ ), .A3(\EXU/CSRControl/_0431_ ), .ZN(\EXU/CSRControl/_0432_ ) );
INV_X1 \EXU/CSRControl/_2328_ ( .A(\EXU/CSRControl/_0288_ ), .ZN(\EXU/CSRControl/_0433_ ) );
OAI211_X2 \EXU/CSRControl/_2329_ ( .A(\EXU/CSRControl/_0432_ ), .B(\EXU/CSRControl/_1213_ ), .C1(\EXU/CSRControl/_0433_ ), .C2(\EXU/CSRControl/_1215_ ), .ZN(\EXU/CSRControl/_0434_ ) );
OR3_X1 \EXU/CSRControl/_2330_ ( .A1(\EXU/CSRControl/_1273_ ), .A2(\EXU/CSRControl/_0274_ ), .A3(\EXU/CSRControl/_0433_ ), .ZN(\EXU/CSRControl/_0435_ ) );
AND2_X2 \EXU/CSRControl/_2331_ ( .A1(\EXU/CSRControl/_0434_ ), .A2(\EXU/CSRControl/_0435_ ), .ZN(\EXU/CSRControl/_0436_ ) );
AOI21_X1 \EXU/CSRControl/_2332_ ( .A(\EXU/CSRControl/_0427_ ), .B1(\EXU/CSRControl/_0436_ ), .B2(\EXU/CSRControl/_1276_ ), .ZN(\EXU/CSRControl/_0025_ ) );
AOI22_X1 \EXU/CSRControl/_2333_ ( .A1(\EXU/CSRControl/_1278_ ), .A2(\EXU/CSRControl/_0210_ ), .B1(\EXU/CSRControl/_1183_ ), .B2(\EXU/CSRControl/_0242_ ), .ZN(\EXU/CSRControl/_0437_ ) );
AOI22_X1 \EXU/CSRControl/_2334_ ( .A1(\EXU/CSRControl/_1205_ ), .A2(\EXU/CSRControl/_0146_ ), .B1(\EXU/CSRControl/_1191_ ), .B2(\EXU/CSRControl/_1147_ ), .ZN(\EXU/CSRControl/_0438_ ) );
NAND3_X1 \EXU/CSRControl/_2335_ ( .A1(\EXU/CSRControl/_1234_ ), .A2(\EXU/CSRControl/_0178_ ), .A3(\EXU/CSRControl/_1235_ ), .ZN(\EXU/CSRControl/_0439_ ) );
NAND3_X1 \EXU/CSRControl/_2336_ ( .A1(\EXU/CSRControl/_0437_ ), .A2(\EXU/CSRControl/_0438_ ), .A3(\EXU/CSRControl/_0439_ ), .ZN(\EXU/CSRControl/_0440_ ) );
NAND3_X1 \EXU/CSRControl/_2337_ ( .A1(\EXU/CSRControl/_0800_ ), .A2(\EXU/CSRControl/_0272_ ), .A3(\EXU/CSRControl/_0289_ ), .ZN(\EXU/CSRControl/_0441_ ) );
NAND3_X1 \EXU/CSRControl/_2338_ ( .A1(\EXU/CSRControl/_0440_ ), .A2(\EXU/CSRControl/_1213_ ), .A3(\EXU/CSRControl/_0441_ ), .ZN(\EXU/CSRControl/_0442_ ) );
NAND2_X1 \EXU/CSRControl/_2339_ ( .A1(\EXU/CSRControl/_1244_ ), .A2(\EXU/CSRControl/_0289_ ), .ZN(\EXU/CSRControl/_0443_ ) );
AND3_X1 \EXU/CSRControl/_2340_ ( .A1(\EXU/CSRControl/_0442_ ), .A2(\EXU/CSRControl/_1243_ ), .A3(\EXU/CSRControl/_0443_ ), .ZN(\EXU/CSRControl/_0444_ ) );
OAI21_X1 \EXU/CSRControl/_2341_ ( .A(\EXU/CSRControl/_1223_ ), .B1(\EXU/CSRControl/_1247_ ), .B2(\EXU/CSRControl/_0242_ ), .ZN(\EXU/CSRControl/_0445_ ) );
NOR2_X1 \EXU/CSRControl/_2342_ ( .A1(\EXU/CSRControl/_0444_ ), .A2(\EXU/CSRControl/_0445_ ), .ZN(\EXU/CSRControl/_0026_ ) );
INV_X1 \EXU/CSRControl/_2343_ ( .A(\EXU/CSRControl/_0290_ ), .ZN(\EXU/CSRControl/_0446_ ) );
NAND2_X1 \EXU/CSRControl/_2344_ ( .A1(\EXU/CSRControl/_1231_ ), .A2(\EXU/CSRControl/_0243_ ), .ZN(\EXU/CSRControl/_0447_ ) );
NAND3_X1 \EXU/CSRControl/_2345_ ( .A1(\EXU/CSRControl/_1234_ ), .A2(\EXU/CSRControl/_0179_ ), .A3(\EXU/CSRControl/_1235_ ), .ZN(\EXU/CSRControl/_0448_ ) );
NAND2_X1 \EXU/CSRControl/_2346_ ( .A1(\EXU/CSRControl/_0447_ ), .A2(\EXU/CSRControl/_0448_ ), .ZN(\EXU/CSRControl/_0449_ ) );
NAND3_X1 \EXU/CSRControl/_2347_ ( .A1(\EXU/CSRControl/_1228_ ), .A2(\EXU/CSRControl/_1229_ ), .A3(\EXU/CSRControl/_0147_ ), .ZN(\EXU/CSRControl/_0450_ ) );
NAND3_X1 \EXU/CSRControl/_2348_ ( .A1(\EXU/CSRControl/_1237_ ), .A2(\EXU/CSRControl/_1269_ ), .A3(\EXU/CSRControl/_0211_ ), .ZN(\EXU/CSRControl/_0451_ ) );
NAND2_X1 \EXU/CSRControl/_2349_ ( .A1(\EXU/CSRControl/_0450_ ), .A2(\EXU/CSRControl/_0451_ ), .ZN(\EXU/CSRControl/_0452_ ) );
OAI221_X1 \EXU/CSRControl/_2350_ ( .A(\EXU/CSRControl/_1263_ ), .B1(\EXU/CSRControl/_0446_ ), .B2(\EXU/CSRControl/_1215_ ), .C1(\EXU/CSRControl/_0449_ ), .C2(\EXU/CSRControl/_0452_ ), .ZN(\EXU/CSRControl/_0453_ ) );
OR3_X1 \EXU/CSRControl/_2351_ ( .A1(\EXU/CSRControl/_1273_ ), .A2(\EXU/CSRControl/_0274_ ), .A3(\EXU/CSRControl/_0446_ ), .ZN(\EXU/CSRControl/_0454_ ) );
AND3_X1 \EXU/CSRControl/_2352_ ( .A1(\EXU/CSRControl/_0453_ ), .A2(\EXU/CSRControl/_1243_ ), .A3(\EXU/CSRControl/_0454_ ), .ZN(\EXU/CSRControl/_0455_ ) );
OAI21_X1 \EXU/CSRControl/_2353_ ( .A(\EXU/CSRControl/_1223_ ), .B1(\EXU/CSRControl/_1247_ ), .B2(\EXU/CSRControl/_0243_ ), .ZN(\EXU/CSRControl/_0456_ ) );
NOR2_X1 \EXU/CSRControl/_2354_ ( .A1(\EXU/CSRControl/_0455_ ), .A2(\EXU/CSRControl/_0456_ ), .ZN(\EXU/CSRControl/_0027_ ) );
BUF_X4 \EXU/CSRControl/_2355_ ( .A(\EXU/CSRControl/_1221_ ), .Z(\EXU/CSRControl/_0457_ ) );
OAI21_X1 \EXU/CSRControl/_2356_ ( .A(\EXU/CSRControl/_0457_ ), .B1(\EXU/CSRControl/_1261_ ), .B2(\EXU/CSRControl/_0244_ ), .ZN(\EXU/CSRControl/_0458_ ) );
AOI22_X1 \EXU/CSRControl/_2357_ ( .A1(\EXU/CSRControl/_1205_ ), .A2(\EXU/CSRControl/_0148_ ), .B1(\EXU/CSRControl/_1139_ ), .B2(\EXU/CSRControl/_0244_ ), .ZN(\EXU/CSRControl/_0459_ ) );
AND3_X1 \EXU/CSRControl/_2358_ ( .A1(\EXU/CSRControl/_1207_ ), .A2(\EXU/CSRControl/_1208_ ), .A3(\EXU/CSRControl/_0212_ ), .ZN(\EXU/CSRControl/_0460_ ) );
NOR2_X1 \EXU/CSRControl/_2359_ ( .A1(\EXU/CSRControl/_0460_ ), .A2(\EXU/CSRControl/_1148_ ), .ZN(\EXU/CSRControl/_0461_ ) );
NAND3_X1 \EXU/CSRControl/_2360_ ( .A1(\EXU/CSRControl/_1187_ ), .A2(\EXU/CSRControl/_0180_ ), .A3(\EXU/CSRControl/_1189_ ), .ZN(\EXU/CSRControl/_0462_ ) );
NAND3_X1 \EXU/CSRControl/_2361_ ( .A1(\EXU/CSRControl/_0459_ ), .A2(\EXU/CSRControl/_0461_ ), .A3(\EXU/CSRControl/_0462_ ), .ZN(\EXU/CSRControl/_0463_ ) );
INV_X1 \EXU/CSRControl/_2362_ ( .A(\EXU/CSRControl/_0291_ ), .ZN(\EXU/CSRControl/_0464_ ) );
OAI211_X2 \EXU/CSRControl/_2363_ ( .A(\EXU/CSRControl/_0463_ ), .B(\EXU/CSRControl/_1263_ ), .C1(\EXU/CSRControl/_0464_ ), .C2(\EXU/CSRControl/_1215_ ), .ZN(\EXU/CSRControl/_0465_ ) );
OR3_X1 \EXU/CSRControl/_2364_ ( .A1(\EXU/CSRControl/_1174_ ), .A2(\EXU/CSRControl/_0274_ ), .A3(\EXU/CSRControl/_0464_ ), .ZN(\EXU/CSRControl/_0466_ ) );
AND2_X2 \EXU/CSRControl/_2365_ ( .A1(\EXU/CSRControl/_0465_ ), .A2(\EXU/CSRControl/_0466_ ), .ZN(\EXU/CSRControl/_0467_ ) );
AOI21_X1 \EXU/CSRControl/_2366_ ( .A(\EXU/CSRControl/_0458_ ), .B1(\EXU/CSRControl/_0467_ ), .B2(\EXU/CSRControl/_1276_ ), .ZN(\EXU/CSRControl/_0028_ ) );
NAND3_X1 \EXU/CSRControl/_2367_ ( .A1(\EXU/CSRControl/_0799_ ), .A2(\EXU/CSRControl/_0272_ ), .A3(\EXU/CSRControl/_0292_ ), .ZN(\EXU/CSRControl/_0468_ ) );
NAND2_X1 \EXU/CSRControl/_2368_ ( .A1(\EXU/CSRControl/_1231_ ), .A2(\EXU/CSRControl/_0245_ ), .ZN(\EXU/CSRControl/_0469_ ) );
NAND3_X1 \EXU/CSRControl/_2369_ ( .A1(\EXU/CSRControl/_1234_ ), .A2(\EXU/CSRControl/_0181_ ), .A3(\EXU/CSRControl/_1235_ ), .ZN(\EXU/CSRControl/_0470_ ) );
NAND2_X1 \EXU/CSRControl/_2370_ ( .A1(\EXU/CSRControl/_0469_ ), .A2(\EXU/CSRControl/_0470_ ), .ZN(\EXU/CSRControl/_0471_ ) );
NAND3_X1 \EXU/CSRControl/_2371_ ( .A1(\EXU/CSRControl/_1228_ ), .A2(\EXU/CSRControl/_1229_ ), .A3(\EXU/CSRControl/_0149_ ), .ZN(\EXU/CSRControl/_0472_ ) );
NAND3_X1 \EXU/CSRControl/_2372_ ( .A1(\EXU/CSRControl/_1237_ ), .A2(\EXU/CSRControl/_1229_ ), .A3(\EXU/CSRControl/_0213_ ), .ZN(\EXU/CSRControl/_0473_ ) );
NAND2_X1 \EXU/CSRControl/_2373_ ( .A1(\EXU/CSRControl/_0472_ ), .A2(\EXU/CSRControl/_0473_ ), .ZN(\EXU/CSRControl/_0474_ ) );
OAI211_X2 \EXU/CSRControl/_2374_ ( .A(\EXU/CSRControl/_1213_ ), .B(\EXU/CSRControl/_0468_ ), .C1(\EXU/CSRControl/_0471_ ), .C2(\EXU/CSRControl/_0474_ ), .ZN(\EXU/CSRControl/_0475_ ) );
NAND2_X1 \EXU/CSRControl/_2375_ ( .A1(\EXU/CSRControl/_1244_ ), .A2(\EXU/CSRControl/_0292_ ), .ZN(\EXU/CSRControl/_0476_ ) );
AND3_X1 \EXU/CSRControl/_2376_ ( .A1(\EXU/CSRControl/_0475_ ), .A2(\EXU/CSRControl/_1243_ ), .A3(\EXU/CSRControl/_0476_ ), .ZN(\EXU/CSRControl/_0477_ ) );
OAI21_X1 \EXU/CSRControl/_2377_ ( .A(\EXU/CSRControl/_1223_ ), .B1(\EXU/CSRControl/_1247_ ), .B2(\EXU/CSRControl/_0245_ ), .ZN(\EXU/CSRControl/_0478_ ) );
NOR2_X1 \EXU/CSRControl/_2378_ ( .A1(\EXU/CSRControl/_0477_ ), .A2(\EXU/CSRControl/_0478_ ), .ZN(\EXU/CSRControl/_0029_ ) );
NAND3_X1 \EXU/CSRControl/_2379_ ( .A1(\EXU/CSRControl/_0799_ ), .A2(\EXU/CSRControl/_0272_ ), .A3(\EXU/CSRControl/_0293_ ), .ZN(\EXU/CSRControl/_0479_ ) );
INV_X1 \EXU/CSRControl/_2380_ ( .A(\EXU/CSRControl/_0246_ ), .ZN(\EXU/CSRControl/_0480_ ) );
OR3_X1 \EXU/CSRControl/_2381_ ( .A1(\EXU/CSRControl/_1137_ ), .A2(\EXU/CSRControl/_0480_ ), .A3(\EXU/CSRControl/_1138_ ), .ZN(\EXU/CSRControl/_0481_ ) );
NAND3_X1 \EXU/CSRControl/_2382_ ( .A1(\EXU/CSRControl/_1186_ ), .A2(\EXU/CSRControl/_0182_ ), .A3(\EXU/CSRControl/_1188_ ), .ZN(\EXU/CSRControl/_0482_ ) );
NAND2_X1 \EXU/CSRControl/_2383_ ( .A1(\EXU/CSRControl/_0481_ ), .A2(\EXU/CSRControl/_0482_ ), .ZN(\EXU/CSRControl/_0483_ ) );
NAND3_X1 \EXU/CSRControl/_2384_ ( .A1(\EXU/CSRControl/_1193_ ), .A2(\EXU/CSRControl/_0874_ ), .A3(\EXU/CSRControl/_0150_ ), .ZN(\EXU/CSRControl/_0484_ ) );
NAND3_X1 \EXU/CSRControl/_2385_ ( .A1(\EXU/CSRControl/_1191_ ), .A2(\EXU/CSRControl/_1117_ ), .A3(\EXU/CSRControl/_0214_ ), .ZN(\EXU/CSRControl/_0485_ ) );
NAND2_X1 \EXU/CSRControl/_2386_ ( .A1(\EXU/CSRControl/_0484_ ), .A2(\EXU/CSRControl/_0485_ ), .ZN(\EXU/CSRControl/_0486_ ) );
OAI211_X2 \EXU/CSRControl/_2387_ ( .A(\EXU/CSRControl/_1181_ ), .B(\EXU/CSRControl/_0479_ ), .C1(\EXU/CSRControl/_0483_ ), .C2(\EXU/CSRControl/_0486_ ), .ZN(\EXU/CSRControl/_0487_ ) );
NAND2_X1 \EXU/CSRControl/_2388_ ( .A1(\EXU/CSRControl/_1155_ ), .A2(\EXU/CSRControl/_0293_ ), .ZN(\EXU/CSRControl/_0488_ ) );
AND3_X1 \EXU/CSRControl/_2389_ ( .A1(\EXU/CSRControl/_0487_ ), .A2(\EXU/CSRControl/_1241_ ), .A3(\EXU/CSRControl/_0488_ ), .ZN(\EXU/CSRControl/_0489_ ) );
AOI211_X2 \EXU/CSRControl/_2390_ ( .A(\EXU/CSRControl/_1374_ ), .B(\EXU/CSRControl/_0489_ ), .C1(\EXU/CSRControl/_0480_ ), .C2(\EXU/CSRControl/_1203_ ), .ZN(\EXU/CSRControl/_0030_ ) );
INV_X1 \EXU/CSRControl/_2391_ ( .A(\EXU/CSRControl/_0294_ ), .ZN(\EXU/CSRControl/_0490_ ) );
NAND2_X1 \EXU/CSRControl/_2392_ ( .A1(\EXU/CSRControl/_1231_ ), .A2(\EXU/CSRControl/_0247_ ), .ZN(\EXU/CSRControl/_0491_ ) );
NAND3_X1 \EXU/CSRControl/_2393_ ( .A1(\EXU/CSRControl/_1237_ ), .A2(\EXU/CSRControl/_1269_ ), .A3(\EXU/CSRControl/_0215_ ), .ZN(\EXU/CSRControl/_0492_ ) );
NAND3_X1 \EXU/CSRControl/_2394_ ( .A1(\EXU/CSRControl/_1228_ ), .A2(\EXU/CSRControl/_1269_ ), .A3(\EXU/CSRControl/_0151_ ), .ZN(\EXU/CSRControl/_0493_ ) );
NAND3_X1 \EXU/CSRControl/_2395_ ( .A1(\EXU/CSRControl/_0491_ ), .A2(\EXU/CSRControl/_0492_ ), .A3(\EXU/CSRControl/_0493_ ), .ZN(\EXU/CSRControl/_0494_ ) );
NAND3_X1 \EXU/CSRControl/_2396_ ( .A1(\EXU/CSRControl/_1187_ ), .A2(\EXU/CSRControl/_0183_ ), .A3(\EXU/CSRControl/_1189_ ), .ZN(\EXU/CSRControl/_0495_ ) );
NAND2_X1 \EXU/CSRControl/_2397_ ( .A1(\EXU/CSRControl/_1149_ ), .A2(\EXU/CSRControl/_0495_ ), .ZN(\EXU/CSRControl/_0496_ ) );
OAI221_X1 \EXU/CSRControl/_2398_ ( .A(\EXU/CSRControl/_1263_ ), .B1(\EXU/CSRControl/_0490_ ), .B2(\EXU/CSRControl/_1215_ ), .C1(\EXU/CSRControl/_0494_ ), .C2(\EXU/CSRControl/_0496_ ), .ZN(\EXU/CSRControl/_0497_ ) );
OR3_X1 \EXU/CSRControl/_2399_ ( .A1(\EXU/CSRControl/_1273_ ), .A2(\EXU/CSRControl/_0274_ ), .A3(\EXU/CSRControl/_0490_ ), .ZN(\EXU/CSRControl/_0498_ ) );
AND3_X1 \EXU/CSRControl/_2400_ ( .A1(\EXU/CSRControl/_0497_ ), .A2(\EXU/CSRControl/_1243_ ), .A3(\EXU/CSRControl/_0498_ ), .ZN(\EXU/CSRControl/_0499_ ) );
OAI21_X1 \EXU/CSRControl/_2401_ ( .A(\EXU/CSRControl/_1223_ ), .B1(\EXU/CSRControl/_1247_ ), .B2(\EXU/CSRControl/_0247_ ), .ZN(\EXU/CSRControl/_0500_ ) );
NOR2_X1 \EXU/CSRControl/_2402_ ( .A1(\EXU/CSRControl/_0499_ ), .A2(\EXU/CSRControl/_0500_ ), .ZN(\EXU/CSRControl/_0031_ ) );
AOI22_X1 \EXU/CSRControl/_2403_ ( .A1(\EXU/CSRControl/_1205_ ), .A2(\EXU/CSRControl/_0152_ ), .B1(\EXU/CSRControl/_1183_ ), .B2(\EXU/CSRControl/_0248_ ), .ZN(\EXU/CSRControl/_0501_ ) );
AND3_X1 \EXU/CSRControl/_2404_ ( .A1(\EXU/CSRControl/_1207_ ), .A2(\EXU/CSRControl/_1208_ ), .A3(\EXU/CSRControl/_0216_ ), .ZN(\EXU/CSRControl/_0502_ ) );
NOR2_X1 \EXU/CSRControl/_2405_ ( .A1(\EXU/CSRControl/_0502_ ), .A2(\EXU/CSRControl/_1148_ ), .ZN(\EXU/CSRControl/_0503_ ) );
NAND3_X1 \EXU/CSRControl/_2406_ ( .A1(\EXU/CSRControl/_1234_ ), .A2(\EXU/CSRControl/_0184_ ), .A3(\EXU/CSRControl/_1235_ ), .ZN(\EXU/CSRControl/_0504_ ) );
NAND3_X1 \EXU/CSRControl/_2407_ ( .A1(\EXU/CSRControl/_0501_ ), .A2(\EXU/CSRControl/_0503_ ), .A3(\EXU/CSRControl/_0504_ ), .ZN(\EXU/CSRControl/_0505_ ) );
NAND3_X1 \EXU/CSRControl/_2408_ ( .A1(\EXU/CSRControl/_0800_ ), .A2(\EXU/CSRControl/_0272_ ), .A3(\EXU/CSRControl/_0295_ ), .ZN(\EXU/CSRControl/_0506_ ) );
NAND3_X1 \EXU/CSRControl/_2409_ ( .A1(\EXU/CSRControl/_0505_ ), .A2(\EXU/CSRControl/_1213_ ), .A3(\EXU/CSRControl/_0506_ ), .ZN(\EXU/CSRControl/_0507_ ) );
NAND2_X1 \EXU/CSRControl/_2410_ ( .A1(\EXU/CSRControl/_1244_ ), .A2(\EXU/CSRControl/_0295_ ), .ZN(\EXU/CSRControl/_0508_ ) );
AND3_X1 \EXU/CSRControl/_2411_ ( .A1(\EXU/CSRControl/_0507_ ), .A2(\EXU/CSRControl/_1242_ ), .A3(\EXU/CSRControl/_0508_ ), .ZN(\EXU/CSRControl/_0509_ ) );
OAI21_X1 \EXU/CSRControl/_2412_ ( .A(\EXU/CSRControl/_1223_ ), .B1(\EXU/CSRControl/_1247_ ), .B2(\EXU/CSRControl/_0248_ ), .ZN(\EXU/CSRControl/_0510_ ) );
NOR2_X1 \EXU/CSRControl/_2413_ ( .A1(\EXU/CSRControl/_0509_ ), .A2(\EXU/CSRControl/_0510_ ), .ZN(\EXU/CSRControl/_0032_ ) );
OAI21_X1 \EXU/CSRControl/_2414_ ( .A(\EXU/CSRControl/_0457_ ), .B1(\EXU/CSRControl/_1243_ ), .B2(\EXU/CSRControl/_0249_ ), .ZN(\EXU/CSRControl/_0511_ ) );
AOI22_X1 \EXU/CSRControl/_2415_ ( .A1(\EXU/CSRControl/_1205_ ), .A2(\EXU/CSRControl/_0153_ ), .B1(\EXU/CSRControl/_1139_ ), .B2(\EXU/CSRControl/_0249_ ), .ZN(\EXU/CSRControl/_0512_ ) );
AND3_X2 \EXU/CSRControl/_2416_ ( .A1(\EXU/CSRControl/_1207_ ), .A2(\EXU/CSRControl/_1208_ ), .A3(\EXU/CSRControl/_0217_ ), .ZN(\EXU/CSRControl/_0513_ ) );
NOR2_X1 \EXU/CSRControl/_2417_ ( .A1(\EXU/CSRControl/_0513_ ), .A2(\EXU/CSRControl/_1148_ ), .ZN(\EXU/CSRControl/_0514_ ) );
NAND3_X1 \EXU/CSRControl/_2418_ ( .A1(\EXU/CSRControl/_1187_ ), .A2(\EXU/CSRControl/_0185_ ), .A3(\EXU/CSRControl/_1189_ ), .ZN(\EXU/CSRControl/_0515_ ) );
NAND3_X1 \EXU/CSRControl/_2419_ ( .A1(\EXU/CSRControl/_0512_ ), .A2(\EXU/CSRControl/_0514_ ), .A3(\EXU/CSRControl/_0515_ ), .ZN(\EXU/CSRControl/_0516_ ) );
INV_X1 \EXU/CSRControl/_2420_ ( .A(\EXU/CSRControl/_0296_ ), .ZN(\EXU/CSRControl/_0517_ ) );
OAI211_X2 \EXU/CSRControl/_2421_ ( .A(\EXU/CSRControl/_0516_ ), .B(\EXU/CSRControl/_1263_ ), .C1(\EXU/CSRControl/_0517_ ), .C2(\EXU/CSRControl/_1215_ ), .ZN(\EXU/CSRControl/_0518_ ) );
OR3_X1 \EXU/CSRControl/_2422_ ( .A1(\EXU/CSRControl/_1174_ ), .A2(\EXU/CSRControl/_0274_ ), .A3(\EXU/CSRControl/_0517_ ), .ZN(\EXU/CSRControl/_0519_ ) );
AND2_X2 \EXU/CSRControl/_2423_ ( .A1(\EXU/CSRControl/_0518_ ), .A2(\EXU/CSRControl/_0519_ ), .ZN(\EXU/CSRControl/_0520_ ) );
AOI21_X1 \EXU/CSRControl/_2424_ ( .A(\EXU/CSRControl/_0511_ ), .B1(\EXU/CSRControl/_0520_ ), .B2(\EXU/CSRControl/_1247_ ), .ZN(\EXU/CSRControl/_0033_ ) );
OAI21_X1 \EXU/CSRControl/_2425_ ( .A(\EXU/CSRControl/_0457_ ), .B1(\EXU/CSRControl/_1243_ ), .B2(\EXU/CSRControl/_0251_ ), .ZN(\EXU/CSRControl/_0521_ ) );
AOI22_X1 \EXU/CSRControl/_2426_ ( .A1(\EXU/CSRControl/_1205_ ), .A2(\EXU/CSRControl/_0155_ ), .B1(\EXU/CSRControl/_1183_ ), .B2(\EXU/CSRControl/_0251_ ), .ZN(\EXU/CSRControl/_0522_ ) );
AND3_X1 \EXU/CSRControl/_2427_ ( .A1(\EXU/CSRControl/_1207_ ), .A2(\EXU/CSRControl/_1208_ ), .A3(\EXU/CSRControl/_0219_ ), .ZN(\EXU/CSRControl/_0523_ ) );
NOR2_X1 \EXU/CSRControl/_2428_ ( .A1(\EXU/CSRControl/_0523_ ), .A2(\EXU/CSRControl/_1148_ ), .ZN(\EXU/CSRControl/_0524_ ) );
NAND3_X1 \EXU/CSRControl/_2429_ ( .A1(\EXU/CSRControl/_1234_ ), .A2(\EXU/CSRControl/_0187_ ), .A3(\EXU/CSRControl/_1235_ ), .ZN(\EXU/CSRControl/_0525_ ) );
NAND3_X1 \EXU/CSRControl/_2430_ ( .A1(\EXU/CSRControl/_0522_ ), .A2(\EXU/CSRControl/_0524_ ), .A3(\EXU/CSRControl/_0525_ ), .ZN(\EXU/CSRControl/_0526_ ) );
NAND3_X1 \EXU/CSRControl/_2431_ ( .A1(\EXU/CSRControl/_0799_ ), .A2(\EXU/CSRControl/_0272_ ), .A3(\EXU/CSRControl/_0298_ ), .ZN(\EXU/CSRControl/_0527_ ) );
NAND3_X1 \EXU/CSRControl/_2432_ ( .A1(\EXU/CSRControl/_0526_ ), .A2(\EXU/CSRControl/_1213_ ), .A3(\EXU/CSRControl/_0527_ ), .ZN(\EXU/CSRControl/_0528_ ) );
NAND2_X1 \EXU/CSRControl/_2433_ ( .A1(\EXU/CSRControl/_1244_ ), .A2(\EXU/CSRControl/_0298_ ), .ZN(\EXU/CSRControl/_0529_ ) );
AND2_X1 \EXU/CSRControl/_2434_ ( .A1(\EXU/CSRControl/_0528_ ), .A2(\EXU/CSRControl/_0529_ ), .ZN(\EXU/CSRControl/_0530_ ) );
AOI21_X1 \EXU/CSRControl/_2435_ ( .A(\EXU/CSRControl/_0521_ ), .B1(\EXU/CSRControl/_0530_ ), .B2(\EXU/CSRControl/_1247_ ), .ZN(\EXU/CSRControl/_0034_ ) );
INV_X1 \EXU/CSRControl/_2436_ ( .A(\EXU/CSRControl/_0299_ ), .ZN(\EXU/CSRControl/_0531_ ) );
INV_X1 \EXU/CSRControl/_2437_ ( .A(\EXU/CSRControl/_0252_ ), .ZN(\EXU/CSRControl/_0532_ ) );
OR3_X1 \EXU/CSRControl/_2438_ ( .A1(\EXU/CSRControl/_1137_ ), .A2(\EXU/CSRControl/_0532_ ), .A3(\EXU/CSRControl/_1138_ ), .ZN(\EXU/CSRControl/_0533_ ) );
NAND3_X1 \EXU/CSRControl/_2439_ ( .A1(\EXU/CSRControl/_1193_ ), .A2(\EXU/CSRControl/_0874_ ), .A3(\EXU/CSRControl/_0156_ ), .ZN(\EXU/CSRControl/_0534_ ) );
NAND2_X1 \EXU/CSRControl/_2440_ ( .A1(\EXU/CSRControl/_0533_ ), .A2(\EXU/CSRControl/_0534_ ), .ZN(\EXU/CSRControl/_0535_ ) );
NAND3_X1 \EXU/CSRControl/_2441_ ( .A1(\EXU/CSRControl/_1186_ ), .A2(\EXU/CSRControl/_0188_ ), .A3(\EXU/CSRControl/_1188_ ), .ZN(\EXU/CSRControl/_0536_ ) );
NAND3_X1 \EXU/CSRControl/_2442_ ( .A1(\EXU/CSRControl/_1207_ ), .A2(\EXU/CSRControl/_1208_ ), .A3(\EXU/CSRControl/_0220_ ), .ZN(\EXU/CSRControl/_0537_ ) );
NAND2_X1 \EXU/CSRControl/_2443_ ( .A1(\EXU/CSRControl/_0536_ ), .A2(\EXU/CSRControl/_0537_ ), .ZN(\EXU/CSRControl/_0538_ ) );
OAI221_X1 \EXU/CSRControl/_2444_ ( .A(\EXU/CSRControl/_1181_ ), .B1(\EXU/CSRControl/_0531_ ), .B2(\EXU/CSRControl/_1166_ ), .C1(\EXU/CSRControl/_0535_ ), .C2(\EXU/CSRControl/_0538_ ), .ZN(\EXU/CSRControl/_0539_ ) );
OR3_X1 \EXU/CSRControl/_2445_ ( .A1(\EXU/CSRControl/_1174_ ), .A2(\EXU/CSRControl/_0274_ ), .A3(\EXU/CSRControl/_0531_ ), .ZN(\EXU/CSRControl/_0540_ ) );
AND3_X1 \EXU/CSRControl/_2446_ ( .A1(\EXU/CSRControl/_0539_ ), .A2(\EXU/CSRControl/_1241_ ), .A3(\EXU/CSRControl/_0540_ ), .ZN(\EXU/CSRControl/_0541_ ) );
AOI211_X2 \EXU/CSRControl/_2447_ ( .A(\EXU/CSRControl/_1374_ ), .B(\EXU/CSRControl/_0541_ ), .C1(\EXU/CSRControl/_0532_ ), .C2(\EXU/CSRControl/_1203_ ), .ZN(\EXU/CSRControl/_0035_ ) );
BUF_X4 \EXU/CSRControl/_2448_ ( .A(\EXU/CSRControl/_1311_ ), .Z(\EXU/CSRControl/_0542_ ) );
CLKBUF_X2 \EXU/CSRControl/_2449_ ( .A(\EXU/CSRControl/_0542_ ), .Z(\EXU/CSRControl/_0543_ ) );
AND3_X1 \EXU/CSRControl/_2450_ ( .A1(\EXU/CSRControl/_1240_ ), .A2(\EXU/CSRControl/_0543_ ), .A3(\EXU/CSRControl/_1245_ ), .ZN(\EXU/CSRControl/_0544_ ) );
BUF_X4 \EXU/CSRControl/_2451_ ( .A(\EXU/CSRControl/_0542_ ), .Z(\EXU/CSRControl/_0545_ ) );
OAI21_X1 \EXU/CSRControl/_2452_ ( .A(\EXU/CSRControl/_1223_ ), .B1(\EXU/CSRControl/_0545_ ), .B2(\EXU/CSRControl/_0164_ ), .ZN(\EXU/CSRControl/_0546_ ) );
NOR2_X1 \EXU/CSRControl/_2453_ ( .A1(\EXU/CSRControl/_0544_ ), .A2(\EXU/CSRControl/_0546_ ), .ZN(\EXU/CSRControl/_0036_ ) );
AND3_X1 \EXU/CSRControl/_2454_ ( .A1(\EXU/CSRControl/_1257_ ), .A2(\EXU/CSRControl/_0543_ ), .A3(\EXU/CSRControl/_1258_ ), .ZN(\EXU/CSRControl/_0547_ ) );
BUF_X4 \EXU/CSRControl/_2455_ ( .A(\EXU/CSRControl/_1222_ ), .Z(\EXU/CSRControl/_0548_ ) );
OAI21_X1 \EXU/CSRControl/_2456_ ( .A(\EXU/CSRControl/_0548_ ), .B1(\EXU/CSRControl/_0545_ ), .B2(\EXU/CSRControl/_0175_ ), .ZN(\EXU/CSRControl/_0549_ ) );
NOR2_X1 \EXU/CSRControl/_2457_ ( .A1(\EXU/CSRControl/_0547_ ), .A2(\EXU/CSRControl/_0549_ ), .ZN(\EXU/CSRControl/_0037_ ) );
AND3_X1 \EXU/CSRControl/_2458_ ( .A1(\EXU/CSRControl/_1272_ ), .A2(\EXU/CSRControl/_0543_ ), .A3(\EXU/CSRControl/_1274_ ), .ZN(\EXU/CSRControl/_0550_ ) );
OAI21_X1 \EXU/CSRControl/_2459_ ( .A(\EXU/CSRControl/_0548_ ), .B1(\EXU/CSRControl/_0545_ ), .B2(\EXU/CSRControl/_0186_ ), .ZN(\EXU/CSRControl/_0551_ ) );
NOR2_X1 \EXU/CSRControl/_2460_ ( .A1(\EXU/CSRControl/_0550_ ), .A2(\EXU/CSRControl/_0551_ ), .ZN(\EXU/CSRControl/_0038_ ) );
AND3_X1 \EXU/CSRControl/_2461_ ( .A1(\EXU/CSRControl/_1153_ ), .A2(\EXU/CSRControl/_0543_ ), .A3(\EXU/CSRControl/_1156_ ), .ZN(\EXU/CSRControl/_0552_ ) );
OAI21_X1 \EXU/CSRControl/_2462_ ( .A(\EXU/CSRControl/_0548_ ), .B1(\EXU/CSRControl/_0545_ ), .B2(\EXU/CSRControl/_0189_ ), .ZN(\EXU/CSRControl/_0553_ ) );
NOR2_X1 \EXU/CSRControl/_2463_ ( .A1(\EXU/CSRControl/_0552_ ), .A2(\EXU/CSRControl/_0553_ ), .ZN(\EXU/CSRControl/_0039_ ) );
AND3_X1 \EXU/CSRControl/_2464_ ( .A1(\EXU/CSRControl/_1285_ ), .A2(\EXU/CSRControl/_0543_ ), .A3(\EXU/CSRControl/_1286_ ), .ZN(\EXU/CSRControl/_0554_ ) );
OAI21_X1 \EXU/CSRControl/_2465_ ( .A(\EXU/CSRControl/_0548_ ), .B1(\EXU/CSRControl/_0545_ ), .B2(\EXU/CSRControl/_0190_ ), .ZN(\EXU/CSRControl/_0555_ ) );
NOR2_X1 \EXU/CSRControl/_2466_ ( .A1(\EXU/CSRControl/_0554_ ), .A2(\EXU/CSRControl/_0555_ ), .ZN(\EXU/CSRControl/_0040_ ) );
AND3_X1 \EXU/CSRControl/_2467_ ( .A1(\EXU/CSRControl/_1296_ ), .A2(\EXU/CSRControl/_0543_ ), .A3(\EXU/CSRControl/_1297_ ), .ZN(\EXU/CSRControl/_0556_ ) );
OAI21_X1 \EXU/CSRControl/_2468_ ( .A(\EXU/CSRControl/_0548_ ), .B1(\EXU/CSRControl/_0545_ ), .B2(\EXU/CSRControl/_0191_ ), .ZN(\EXU/CSRControl/_0557_ ) );
NOR2_X1 \EXU/CSRControl/_2469_ ( .A1(\EXU/CSRControl/_0556_ ), .A2(\EXU/CSRControl/_0557_ ), .ZN(\EXU/CSRControl/_0041_ ) );
AND3_X1 \EXU/CSRControl/_2470_ ( .A1(\EXU/CSRControl/_1307_ ), .A2(\EXU/CSRControl/_0543_ ), .A3(\EXU/CSRControl/_1308_ ), .ZN(\EXU/CSRControl/_0558_ ) );
OAI21_X1 \EXU/CSRControl/_2471_ ( .A(\EXU/CSRControl/_0548_ ), .B1(\EXU/CSRControl/_0545_ ), .B2(\EXU/CSRControl/_0192_ ), .ZN(\EXU/CSRControl/_0559_ ) );
NOR2_X1 \EXU/CSRControl/_2472_ ( .A1(\EXU/CSRControl/_0558_ ), .A2(\EXU/CSRControl/_0559_ ), .ZN(\EXU/CSRControl/_0042_ ) );
AND3_X1 \EXU/CSRControl/_2473_ ( .A1(\EXU/CSRControl/_1173_ ), .A2(\EXU/CSRControl/_0543_ ), .A3(\EXU/CSRControl/_1175_ ), .ZN(\EXU/CSRControl/_0560_ ) );
OAI21_X1 \EXU/CSRControl/_2474_ ( .A(\EXU/CSRControl/_0548_ ), .B1(\EXU/CSRControl/_0545_ ), .B2(\EXU/CSRControl/_0193_ ), .ZN(\EXU/CSRControl/_0561_ ) );
NOR2_X1 \EXU/CSRControl/_2475_ ( .A1(\EXU/CSRControl/_0560_ ), .A2(\EXU/CSRControl/_0561_ ), .ZN(\EXU/CSRControl/_0043_ ) );
CLKBUF_X2 \EXU/CSRControl/_2476_ ( .A(\EXU/CSRControl/_0542_ ), .Z(\EXU/CSRControl/_0562_ ) );
AND3_X1 \EXU/CSRControl/_2477_ ( .A1(\EXU/CSRControl/_1317_ ), .A2(\EXU/CSRControl/_0562_ ), .A3(\EXU/CSRControl/_1318_ ), .ZN(\EXU/CSRControl/_0563_ ) );
OAI21_X1 \EXU/CSRControl/_2478_ ( .A(\EXU/CSRControl/_0548_ ), .B1(\EXU/CSRControl/_0545_ ), .B2(\EXU/CSRControl/_0194_ ), .ZN(\EXU/CSRControl/_0564_ ) );
NOR2_X1 \EXU/CSRControl/_2479_ ( .A1(\EXU/CSRControl/_0563_ ), .A2(\EXU/CSRControl/_0564_ ), .ZN(\EXU/CSRControl/_0044_ ) );
AND3_X1 \EXU/CSRControl/_2480_ ( .A1(\EXU/CSRControl/_1328_ ), .A2(\EXU/CSRControl/_0562_ ), .A3(\EXU/CSRControl/_1329_ ), .ZN(\EXU/CSRControl/_0565_ ) );
OAI21_X1 \EXU/CSRControl/_2481_ ( .A(\EXU/CSRControl/_0548_ ), .B1(\EXU/CSRControl/_0545_ ), .B2(\EXU/CSRControl/_0195_ ), .ZN(\EXU/CSRControl/_0566_ ) );
NOR2_X1 \EXU/CSRControl/_2482_ ( .A1(\EXU/CSRControl/_0565_ ), .A2(\EXU/CSRControl/_0566_ ), .ZN(\EXU/CSRControl/_0045_ ) );
AND3_X1 \EXU/CSRControl/_2483_ ( .A1(\EXU/CSRControl/_1339_ ), .A2(\EXU/CSRControl/_0562_ ), .A3(\EXU/CSRControl/_1340_ ), .ZN(\EXU/CSRControl/_0567_ ) );
BUF_X4 \EXU/CSRControl/_2484_ ( .A(\EXU/CSRControl/_0542_ ), .Z(\EXU/CSRControl/_0568_ ) );
OAI21_X1 \EXU/CSRControl/_2485_ ( .A(\EXU/CSRControl/_0548_ ), .B1(\EXU/CSRControl/_0568_ ), .B2(\EXU/CSRControl/_0165_ ), .ZN(\EXU/CSRControl/_0569_ ) );
NOR2_X1 \EXU/CSRControl/_2486_ ( .A1(\EXU/CSRControl/_0567_ ), .A2(\EXU/CSRControl/_0569_ ), .ZN(\EXU/CSRControl/_0046_ ) );
AND3_X1 \EXU/CSRControl/_2487_ ( .A1(\EXU/CSRControl/_1196_ ), .A2(\EXU/CSRControl/_0562_ ), .A3(\EXU/CSRControl/_1197_ ), .ZN(\EXU/CSRControl/_0570_ ) );
BUF_X4 \EXU/CSRControl/_2488_ ( .A(\EXU/CSRControl/_1222_ ), .Z(\EXU/CSRControl/_0571_ ) );
OAI21_X1 \EXU/CSRControl/_2489_ ( .A(\EXU/CSRControl/_0571_ ), .B1(\EXU/CSRControl/_0568_ ), .B2(\EXU/CSRControl/_0166_ ), .ZN(\EXU/CSRControl/_0572_ ) );
NOR2_X1 \EXU/CSRControl/_2490_ ( .A1(\EXU/CSRControl/_0570_ ), .A2(\EXU/CSRControl/_0572_ ), .ZN(\EXU/CSRControl/_0047_ ) );
AND3_X1 \EXU/CSRControl/_2491_ ( .A1(\EXU/CSRControl/_1216_ ), .A2(\EXU/CSRControl/_0562_ ), .A3(\EXU/CSRControl/_1217_ ), .ZN(\EXU/CSRControl/_0573_ ) );
OAI21_X1 \EXU/CSRControl/_2492_ ( .A(\EXU/CSRControl/_0571_ ), .B1(\EXU/CSRControl/_0568_ ), .B2(\EXU/CSRControl/_0167_ ), .ZN(\EXU/CSRControl/_0574_ ) );
NOR2_X1 \EXU/CSRControl/_2493_ ( .A1(\EXU/CSRControl/_0573_ ), .A2(\EXU/CSRControl/_0574_ ), .ZN(\EXU/CSRControl/_0048_ ) );
AND3_X1 \EXU/CSRControl/_2494_ ( .A1(\EXU/CSRControl/_1349_ ), .A2(\EXU/CSRControl/_0562_ ), .A3(\EXU/CSRControl/_1350_ ), .ZN(\EXU/CSRControl/_0575_ ) );
OAI21_X1 \EXU/CSRControl/_2495_ ( .A(\EXU/CSRControl/_0571_ ), .B1(\EXU/CSRControl/_0568_ ), .B2(\EXU/CSRControl/_0168_ ), .ZN(\EXU/CSRControl/_0576_ ) );
NOR2_X1 \EXU/CSRControl/_2496_ ( .A1(\EXU/CSRControl/_0575_ ), .A2(\EXU/CSRControl/_0576_ ), .ZN(\EXU/CSRControl/_0049_ ) );
AND3_X1 \EXU/CSRControl/_2497_ ( .A1(\EXU/CSRControl/_1359_ ), .A2(\EXU/CSRControl/_0562_ ), .A3(\EXU/CSRControl/_1360_ ), .ZN(\EXU/CSRControl/_0577_ ) );
OAI21_X1 \EXU/CSRControl/_2498_ ( .A(\EXU/CSRControl/_0571_ ), .B1(\EXU/CSRControl/_0568_ ), .B2(\EXU/CSRControl/_0169_ ), .ZN(\EXU/CSRControl/_0578_ ) );
NOR2_X1 \EXU/CSRControl/_2499_ ( .A1(\EXU/CSRControl/_0577_ ), .A2(\EXU/CSRControl/_0578_ ), .ZN(\EXU/CSRControl/_0050_ ) );
AND3_X1 \EXU/CSRControl/_2500_ ( .A1(\EXU/CSRControl/_1369_ ), .A2(\EXU/CSRControl/_0562_ ), .A3(\EXU/CSRControl/_1370_ ), .ZN(\EXU/CSRControl/_0579_ ) );
OAI21_X1 \EXU/CSRControl/_2501_ ( .A(\EXU/CSRControl/_0571_ ), .B1(\EXU/CSRControl/_0568_ ), .B2(\EXU/CSRControl/_0170_ ), .ZN(\EXU/CSRControl/_0580_ ) );
NOR2_X1 \EXU/CSRControl/_2502_ ( .A1(\EXU/CSRControl/_0579_ ), .A2(\EXU/CSRControl/_0580_ ), .ZN(\EXU/CSRControl/_0051_ ) );
AND3_X1 \EXU/CSRControl/_2503_ ( .A1(\EXU/CSRControl/_0380_ ), .A2(\EXU/CSRControl/_0562_ ), .A3(\EXU/CSRControl/_0381_ ), .ZN(\EXU/CSRControl/_0581_ ) );
OAI21_X1 \EXU/CSRControl/_2504_ ( .A(\EXU/CSRControl/_0571_ ), .B1(\EXU/CSRControl/_0568_ ), .B2(\EXU/CSRControl/_0171_ ), .ZN(\EXU/CSRControl/_0582_ ) );
NOR2_X1 \EXU/CSRControl/_2505_ ( .A1(\EXU/CSRControl/_0581_ ), .A2(\EXU/CSRControl/_0582_ ), .ZN(\EXU/CSRControl/_0052_ ) );
AND3_X1 \EXU/CSRControl/_2506_ ( .A1(\EXU/CSRControl/_0391_ ), .A2(\EXU/CSRControl/_0562_ ), .A3(\EXU/CSRControl/_0392_ ), .ZN(\EXU/CSRControl/_0583_ ) );
OAI21_X1 \EXU/CSRControl/_2507_ ( .A(\EXU/CSRControl/_0571_ ), .B1(\EXU/CSRControl/_0568_ ), .B2(\EXU/CSRControl/_0172_ ), .ZN(\EXU/CSRControl/_0584_ ) );
NOR2_X1 \EXU/CSRControl/_2508_ ( .A1(\EXU/CSRControl/_0583_ ), .A2(\EXU/CSRControl/_0584_ ), .ZN(\EXU/CSRControl/_0053_ ) );
CLKBUF_X2 \EXU/CSRControl/_2509_ ( .A(\EXU/CSRControl/_0542_ ), .Z(\EXU/CSRControl/_0585_ ) );
AND3_X1 \EXU/CSRControl/_2510_ ( .A1(\EXU/CSRControl/_0402_ ), .A2(\EXU/CSRControl/_0585_ ), .A3(\EXU/CSRControl/_0403_ ), .ZN(\EXU/CSRControl/_0586_ ) );
OAI21_X1 \EXU/CSRControl/_2511_ ( .A(\EXU/CSRControl/_0571_ ), .B1(\EXU/CSRControl/_0568_ ), .B2(\EXU/CSRControl/_0173_ ), .ZN(\EXU/CSRControl/_0587_ ) );
NOR2_X1 \EXU/CSRControl/_2512_ ( .A1(\EXU/CSRControl/_0586_ ), .A2(\EXU/CSRControl/_0587_ ), .ZN(\EXU/CSRControl/_0054_ ) );
AND3_X1 \EXU/CSRControl/_2513_ ( .A1(\EXU/CSRControl/_0413_ ), .A2(\EXU/CSRControl/_0585_ ), .A3(\EXU/CSRControl/_0414_ ), .ZN(\EXU/CSRControl/_0588_ ) );
OAI21_X1 \EXU/CSRControl/_2514_ ( .A(\EXU/CSRControl/_0571_ ), .B1(\EXU/CSRControl/_0568_ ), .B2(\EXU/CSRControl/_0174_ ), .ZN(\EXU/CSRControl/_0589_ ) );
NOR2_X1 \EXU/CSRControl/_2515_ ( .A1(\EXU/CSRControl/_0588_ ), .A2(\EXU/CSRControl/_0589_ ), .ZN(\EXU/CSRControl/_0055_ ) );
AND3_X1 \EXU/CSRControl/_2516_ ( .A1(\EXU/CSRControl/_0424_ ), .A2(\EXU/CSRControl/_0585_ ), .A3(\EXU/CSRControl/_0425_ ), .ZN(\EXU/CSRControl/_0590_ ) );
BUF_X4 \EXU/CSRControl/_2517_ ( .A(\EXU/CSRControl/_0542_ ), .Z(\EXU/CSRControl/_0591_ ) );
OAI21_X1 \EXU/CSRControl/_2518_ ( .A(\EXU/CSRControl/_0571_ ), .B1(\EXU/CSRControl/_0591_ ), .B2(\EXU/CSRControl/_0176_ ), .ZN(\EXU/CSRControl/_0592_ ) );
NOR2_X1 \EXU/CSRControl/_2519_ ( .A1(\EXU/CSRControl/_0590_ ), .A2(\EXU/CSRControl/_0592_ ), .ZN(\EXU/CSRControl/_0056_ ) );
AND3_X1 \EXU/CSRControl/_2520_ ( .A1(\EXU/CSRControl/_0434_ ), .A2(\EXU/CSRControl/_0585_ ), .A3(\EXU/CSRControl/_0435_ ), .ZN(\EXU/CSRControl/_0593_ ) );
BUF_X4 \EXU/CSRControl/_2521_ ( .A(\EXU/CSRControl/_1221_ ), .Z(\EXU/CSRControl/_0594_ ) );
OAI21_X1 \EXU/CSRControl/_2522_ ( .A(\EXU/CSRControl/_0594_ ), .B1(\EXU/CSRControl/_0591_ ), .B2(\EXU/CSRControl/_0177_ ), .ZN(\EXU/CSRControl/_0595_ ) );
NOR2_X1 \EXU/CSRControl/_2523_ ( .A1(\EXU/CSRControl/_0593_ ), .A2(\EXU/CSRControl/_0595_ ), .ZN(\EXU/CSRControl/_0057_ ) );
AND3_X1 \EXU/CSRControl/_2524_ ( .A1(\EXU/CSRControl/_0442_ ), .A2(\EXU/CSRControl/_0585_ ), .A3(\EXU/CSRControl/_0443_ ), .ZN(\EXU/CSRControl/_0596_ ) );
OAI21_X1 \EXU/CSRControl/_2525_ ( .A(\EXU/CSRControl/_0594_ ), .B1(\EXU/CSRControl/_0591_ ), .B2(\EXU/CSRControl/_0178_ ), .ZN(\EXU/CSRControl/_0597_ ) );
NOR2_X1 \EXU/CSRControl/_2526_ ( .A1(\EXU/CSRControl/_0596_ ), .A2(\EXU/CSRControl/_0597_ ), .ZN(\EXU/CSRControl/_0058_ ) );
AND3_X1 \EXU/CSRControl/_2527_ ( .A1(\EXU/CSRControl/_0453_ ), .A2(\EXU/CSRControl/_0585_ ), .A3(\EXU/CSRControl/_0454_ ), .ZN(\EXU/CSRControl/_0598_ ) );
OAI21_X1 \EXU/CSRControl/_2528_ ( .A(\EXU/CSRControl/_0594_ ), .B1(\EXU/CSRControl/_0591_ ), .B2(\EXU/CSRControl/_0179_ ), .ZN(\EXU/CSRControl/_0599_ ) );
NOR2_X1 \EXU/CSRControl/_2529_ ( .A1(\EXU/CSRControl/_0598_ ), .A2(\EXU/CSRControl/_0599_ ), .ZN(\EXU/CSRControl/_0059_ ) );
AND3_X1 \EXU/CSRControl/_2530_ ( .A1(\EXU/CSRControl/_0465_ ), .A2(\EXU/CSRControl/_0585_ ), .A3(\EXU/CSRControl/_0466_ ), .ZN(\EXU/CSRControl/_0600_ ) );
OAI21_X1 \EXU/CSRControl/_2531_ ( .A(\EXU/CSRControl/_0594_ ), .B1(\EXU/CSRControl/_0591_ ), .B2(\EXU/CSRControl/_0180_ ), .ZN(\EXU/CSRControl/_0601_ ) );
NOR2_X1 \EXU/CSRControl/_2532_ ( .A1(\EXU/CSRControl/_0600_ ), .A2(\EXU/CSRControl/_0601_ ), .ZN(\EXU/CSRControl/_0060_ ) );
AND3_X1 \EXU/CSRControl/_2533_ ( .A1(\EXU/CSRControl/_0475_ ), .A2(\EXU/CSRControl/_0585_ ), .A3(\EXU/CSRControl/_0476_ ), .ZN(\EXU/CSRControl/_0602_ ) );
OAI21_X1 \EXU/CSRControl/_2534_ ( .A(\EXU/CSRControl/_0594_ ), .B1(\EXU/CSRControl/_0591_ ), .B2(\EXU/CSRControl/_0181_ ), .ZN(\EXU/CSRControl/_0603_ ) );
NOR2_X1 \EXU/CSRControl/_2535_ ( .A1(\EXU/CSRControl/_0602_ ), .A2(\EXU/CSRControl/_0603_ ), .ZN(\EXU/CSRControl/_0061_ ) );
AND3_X1 \EXU/CSRControl/_2536_ ( .A1(\EXU/CSRControl/_0487_ ), .A2(\EXU/CSRControl/_0585_ ), .A3(\EXU/CSRControl/_0488_ ), .ZN(\EXU/CSRControl/_0604_ ) );
OAI21_X1 \EXU/CSRControl/_2537_ ( .A(\EXU/CSRControl/_0594_ ), .B1(\EXU/CSRControl/_0591_ ), .B2(\EXU/CSRControl/_0182_ ), .ZN(\EXU/CSRControl/_0605_ ) );
NOR2_X1 \EXU/CSRControl/_2538_ ( .A1(\EXU/CSRControl/_0604_ ), .A2(\EXU/CSRControl/_0605_ ), .ZN(\EXU/CSRControl/_0062_ ) );
AND3_X1 \EXU/CSRControl/_2539_ ( .A1(\EXU/CSRControl/_0497_ ), .A2(\EXU/CSRControl/_0585_ ), .A3(\EXU/CSRControl/_0498_ ), .ZN(\EXU/CSRControl/_0606_ ) );
OAI21_X1 \EXU/CSRControl/_2540_ ( .A(\EXU/CSRControl/_0594_ ), .B1(\EXU/CSRControl/_0591_ ), .B2(\EXU/CSRControl/_0183_ ), .ZN(\EXU/CSRControl/_0607_ ) );
NOR2_X1 \EXU/CSRControl/_2541_ ( .A1(\EXU/CSRControl/_0606_ ), .A2(\EXU/CSRControl/_0607_ ), .ZN(\EXU/CSRControl/_0063_ ) );
AND3_X1 \EXU/CSRControl/_2542_ ( .A1(\EXU/CSRControl/_0507_ ), .A2(\EXU/CSRControl/_0542_ ), .A3(\EXU/CSRControl/_0508_ ), .ZN(\EXU/CSRControl/_0608_ ) );
OAI21_X1 \EXU/CSRControl/_2543_ ( .A(\EXU/CSRControl/_0594_ ), .B1(\EXU/CSRControl/_0591_ ), .B2(\EXU/CSRControl/_0184_ ), .ZN(\EXU/CSRControl/_0609_ ) );
NOR2_X1 \EXU/CSRControl/_2544_ ( .A1(\EXU/CSRControl/_0608_ ), .A2(\EXU/CSRControl/_0609_ ), .ZN(\EXU/CSRControl/_0064_ ) );
AND3_X1 \EXU/CSRControl/_2545_ ( .A1(\EXU/CSRControl/_0518_ ), .A2(\EXU/CSRControl/_0542_ ), .A3(\EXU/CSRControl/_0519_ ), .ZN(\EXU/CSRControl/_0610_ ) );
OAI21_X1 \EXU/CSRControl/_2546_ ( .A(\EXU/CSRControl/_0594_ ), .B1(\EXU/CSRControl/_0591_ ), .B2(\EXU/CSRControl/_0185_ ), .ZN(\EXU/CSRControl/_0611_ ) );
NOR2_X1 \EXU/CSRControl/_2547_ ( .A1(\EXU/CSRControl/_0610_ ), .A2(\EXU/CSRControl/_0611_ ), .ZN(\EXU/CSRControl/_0065_ ) );
AND3_X1 \EXU/CSRControl/_2548_ ( .A1(\EXU/CSRControl/_0528_ ), .A2(\EXU/CSRControl/_0542_ ), .A3(\EXU/CSRControl/_0529_ ), .ZN(\EXU/CSRControl/_0612_ ) );
OAI21_X1 \EXU/CSRControl/_2549_ ( .A(\EXU/CSRControl/_0594_ ), .B1(\EXU/CSRControl/_0543_ ), .B2(\EXU/CSRControl/_0187_ ), .ZN(\EXU/CSRControl/_0613_ ) );
NOR2_X1 \EXU/CSRControl/_2550_ ( .A1(\EXU/CSRControl/_0612_ ), .A2(\EXU/CSRControl/_0613_ ), .ZN(\EXU/CSRControl/_0066_ ) );
AND3_X1 \EXU/CSRControl/_2551_ ( .A1(\EXU/CSRControl/_0539_ ), .A2(\EXU/CSRControl/_0542_ ), .A3(\EXU/CSRControl/_0540_ ), .ZN(\EXU/CSRControl/_0614_ ) );
OAI21_X1 \EXU/CSRControl/_2552_ ( .A(\EXU/CSRControl/_1260_ ), .B1(\EXU/CSRControl/_0543_ ), .B2(\EXU/CSRControl/_0188_ ), .ZN(\EXU/CSRControl/_0615_ ) );
NOR2_X1 \EXU/CSRControl/_2553_ ( .A1(\EXU/CSRControl/_0614_ ), .A2(\EXU/CSRControl/_0615_ ), .ZN(\EXU/CSRControl/_0067_ ) );
OR2_X1 \EXU/CSRControl/_2554_ ( .A1(\EXU/CSRControl/_1278_ ), .A2(\EXU/CSRControl/_0795_ ), .ZN(\EXU/CSRControl/_0616_ ) );
AOI21_X1 \EXU/CSRControl/_2555_ ( .A(\EXU/CSRControl/_0797_ ), .B1(\EXU/CSRControl/_0272_ ), .B2(\EXU/CSRControl/_0803_ ), .ZN(\EXU/CSRControl/_0617_ ) );
AND2_X2 \EXU/CSRControl/_2556_ ( .A1(\EXU/CSRControl/_0616_ ), .A2(\EXU/CSRControl/_0617_ ), .ZN(\EXU/CSRControl/_0618_ ) );
BUF_X4 \EXU/CSRControl/_2557_ ( .A(\EXU/CSRControl/_0618_ ), .Z(\EXU/CSRControl/_0619_ ) );
OAI21_X1 \EXU/CSRControl/_2558_ ( .A(\EXU/CSRControl/_0457_ ), .B1(\EXU/CSRControl/_0619_ ), .B2(\EXU/CSRControl/_0196_ ), .ZN(\EXU/CSRControl/_0620_ ) );
AND2_X1 \EXU/CSRControl/_2559_ ( .A1(\EXU/CSRControl/_1240_ ), .A2(\EXU/CSRControl/_1245_ ), .ZN(\EXU/CSRControl/_0621_ ) );
OR2_X1 \EXU/CSRControl/_2560_ ( .A1(\EXU/CSRControl/_0621_ ), .A2(\EXU/CSRControl/_1200_ ), .ZN(\EXU/CSRControl/_0622_ ) );
INV_X1 \EXU/CSRControl/_2561_ ( .A(\EXU/CSRControl/_0618_ ), .ZN(\EXU/CSRControl/_0623_ ) );
BUF_X4 \EXU/CSRControl/_2562_ ( .A(\EXU/CSRControl/_0623_ ), .Z(\EXU/CSRControl/_0624_ ) );
BUF_X4 \EXU/CSRControl/_2563_ ( .A(\EXU/CSRControl/_1160_ ), .Z(\EXU/CSRControl/_0625_ ) );
AOI21_X1 \EXU/CSRControl/_2564_ ( .A(\EXU/CSRControl/_0624_ ), .B1(\EXU/CSRControl/_0339_ ), .B2(\EXU/CSRControl/_0625_ ), .ZN(\EXU/CSRControl/_0626_ ) );
AOI21_X1 \EXU/CSRControl/_2565_ ( .A(\EXU/CSRControl/_0620_ ), .B1(\EXU/CSRControl/_0622_ ), .B2(\EXU/CSRControl/_0626_ ), .ZN(\EXU/CSRControl/_0068_ ) );
OAI21_X1 \EXU/CSRControl/_2566_ ( .A(\EXU/CSRControl/_0457_ ), .B1(\EXU/CSRControl/_0619_ ), .B2(\EXU/CSRControl/_0207_ ), .ZN(\EXU/CSRControl/_0627_ ) );
AND2_X1 \EXU/CSRControl/_2567_ ( .A1(\EXU/CSRControl/_1257_ ), .A2(\EXU/CSRControl/_1258_ ), .ZN(\EXU/CSRControl/_0628_ ) );
OR2_X1 \EXU/CSRControl/_2568_ ( .A1(\EXU/CSRControl/_0628_ ), .A2(\EXU/CSRControl/_1200_ ), .ZN(\EXU/CSRControl/_0629_ ) );
AOI21_X1 \EXU/CSRControl/_2569_ ( .A(\EXU/CSRControl/_0624_ ), .B1(\EXU/CSRControl/_0350_ ), .B2(\EXU/CSRControl/_0625_ ), .ZN(\EXU/CSRControl/_0630_ ) );
AOI21_X1 \EXU/CSRControl/_2570_ ( .A(\EXU/CSRControl/_0627_ ), .B1(\EXU/CSRControl/_0629_ ), .B2(\EXU/CSRControl/_0630_ ), .ZN(\EXU/CSRControl/_0069_ ) );
OAI21_X1 \EXU/CSRControl/_2571_ ( .A(\EXU/CSRControl/_0457_ ), .B1(\EXU/CSRControl/_0619_ ), .B2(\EXU/CSRControl/_0218_ ), .ZN(\EXU/CSRControl/_0631_ ) );
OR2_X4 \EXU/CSRControl/_2572_ ( .A1(\EXU/CSRControl/_1275_ ), .A2(\EXU/CSRControl/_1200_ ), .ZN(\EXU/CSRControl/_0632_ ) );
AOI21_X1 \EXU/CSRControl/_2573_ ( .A(\EXU/CSRControl/_0624_ ), .B1(\EXU/CSRControl/_0361_ ), .B2(\EXU/CSRControl/_0625_ ), .ZN(\EXU/CSRControl/_0633_ ) );
AOI21_X1 \EXU/CSRControl/_2574_ ( .A(\EXU/CSRControl/_0631_ ), .B1(\EXU/CSRControl/_0632_ ), .B2(\EXU/CSRControl/_0633_ ), .ZN(\EXU/CSRControl/_0070_ ) );
OAI21_X1 \EXU/CSRControl/_2575_ ( .A(\EXU/CSRControl/_0457_ ), .B1(\EXU/CSRControl/_0619_ ), .B2(\EXU/CSRControl/_0221_ ), .ZN(\EXU/CSRControl/_0634_ ) );
OR2_X1 \EXU/CSRControl/_2576_ ( .A1(\EXU/CSRControl/_1157_ ), .A2(\EXU/CSRControl/_1160_ ), .ZN(\EXU/CSRControl/_0635_ ) );
AOI21_X1 \EXU/CSRControl/_2577_ ( .A(\EXU/CSRControl/_0624_ ), .B1(\EXU/CSRControl/_0364_ ), .B2(\EXU/CSRControl/_0625_ ), .ZN(\EXU/CSRControl/_0636_ ) );
AOI21_X1 \EXU/CSRControl/_2578_ ( .A(\EXU/CSRControl/_0634_ ), .B1(\EXU/CSRControl/_0635_ ), .B2(\EXU/CSRControl/_0636_ ), .ZN(\EXU/CSRControl/_0071_ ) );
OAI21_X1 \EXU/CSRControl/_2579_ ( .A(\EXU/CSRControl/_0457_ ), .B1(\EXU/CSRControl/_0619_ ), .B2(\EXU/CSRControl/_0222_ ), .ZN(\EXU/CSRControl/_0637_ ) );
OR2_X1 \EXU/CSRControl/_2580_ ( .A1(\EXU/CSRControl/_1287_ ), .A2(\EXU/CSRControl/_1200_ ), .ZN(\EXU/CSRControl/_0638_ ) );
AOI21_X1 \EXU/CSRControl/_2581_ ( .A(\EXU/CSRControl/_0624_ ), .B1(\EXU/CSRControl/_0365_ ), .B2(\EXU/CSRControl/_0625_ ), .ZN(\EXU/CSRControl/_0639_ ) );
AOI21_X1 \EXU/CSRControl/_2582_ ( .A(\EXU/CSRControl/_0637_ ), .B1(\EXU/CSRControl/_0638_ ), .B2(\EXU/CSRControl/_0639_ ), .ZN(\EXU/CSRControl/_0072_ ) );
OAI21_X1 \EXU/CSRControl/_2583_ ( .A(\EXU/CSRControl/_0457_ ), .B1(\EXU/CSRControl/_0619_ ), .B2(\EXU/CSRControl/_0223_ ), .ZN(\EXU/CSRControl/_0640_ ) );
OR2_X1 \EXU/CSRControl/_2584_ ( .A1(\EXU/CSRControl/_1298_ ), .A2(\EXU/CSRControl/_1200_ ), .ZN(\EXU/CSRControl/_0641_ ) );
AOI21_X1 \EXU/CSRControl/_2585_ ( .A(\EXU/CSRControl/_0624_ ), .B1(\EXU/CSRControl/_0366_ ), .B2(\EXU/CSRControl/_0625_ ), .ZN(\EXU/CSRControl/_0642_ ) );
AOI21_X1 \EXU/CSRControl/_2586_ ( .A(\EXU/CSRControl/_0640_ ), .B1(\EXU/CSRControl/_0641_ ), .B2(\EXU/CSRControl/_0642_ ), .ZN(\EXU/CSRControl/_0073_ ) );
OAI21_X1 \EXU/CSRControl/_2587_ ( .A(\EXU/CSRControl/_0457_ ), .B1(\EXU/CSRControl/_0619_ ), .B2(\EXU/CSRControl/_0224_ ), .ZN(\EXU/CSRControl/_0643_ ) );
AND2_X1 \EXU/CSRControl/_2588_ ( .A1(\EXU/CSRControl/_1307_ ), .A2(\EXU/CSRControl/_1308_ ), .ZN(\EXU/CSRControl/_0644_ ) );
CLKBUF_X2 \EXU/CSRControl/_2589_ ( .A(\EXU/CSRControl/_0841_ ), .Z(\EXU/CSRControl/_0645_ ) );
OR2_X1 \EXU/CSRControl/_2590_ ( .A1(\EXU/CSRControl/_0644_ ), .A2(\EXU/CSRControl/_0645_ ), .ZN(\EXU/CSRControl/_0646_ ) );
AOI21_X1 \EXU/CSRControl/_2591_ ( .A(\EXU/CSRControl/_0624_ ), .B1(\EXU/CSRControl/_0367_ ), .B2(\EXU/CSRControl/_0625_ ), .ZN(\EXU/CSRControl/_0647_ ) );
AOI21_X1 \EXU/CSRControl/_2592_ ( .A(\EXU/CSRControl/_0643_ ), .B1(\EXU/CSRControl/_0646_ ), .B2(\EXU/CSRControl/_0647_ ), .ZN(\EXU/CSRControl/_0074_ ) );
BUF_X4 \EXU/CSRControl/_2593_ ( .A(\EXU/CSRControl/_1221_ ), .Z(\EXU/CSRControl/_0648_ ) );
OAI21_X1 \EXU/CSRControl/_2594_ ( .A(\EXU/CSRControl/_0648_ ), .B1(\EXU/CSRControl/_0619_ ), .B2(\EXU/CSRControl/_0225_ ), .ZN(\EXU/CSRControl/_0649_ ) );
OR2_X1 \EXU/CSRControl/_2595_ ( .A1(\EXU/CSRControl/_1176_ ), .A2(\EXU/CSRControl/_0645_ ), .ZN(\EXU/CSRControl/_0650_ ) );
AOI21_X1 \EXU/CSRControl/_2596_ ( .A(\EXU/CSRControl/_0624_ ), .B1(\EXU/CSRControl/_0368_ ), .B2(\EXU/CSRControl/_0625_ ), .ZN(\EXU/CSRControl/_0651_ ) );
AOI21_X1 \EXU/CSRControl/_2597_ ( .A(\EXU/CSRControl/_0649_ ), .B1(\EXU/CSRControl/_0650_ ), .B2(\EXU/CSRControl/_0651_ ), .ZN(\EXU/CSRControl/_0075_ ) );
OAI21_X1 \EXU/CSRControl/_2598_ ( .A(\EXU/CSRControl/_0648_ ), .B1(\EXU/CSRControl/_0619_ ), .B2(\EXU/CSRControl/_0226_ ), .ZN(\EXU/CSRControl/_0652_ ) );
OR2_X1 \EXU/CSRControl/_2599_ ( .A1(\EXU/CSRControl/_1319_ ), .A2(\EXU/CSRControl/_0645_ ), .ZN(\EXU/CSRControl/_0653_ ) );
AOI21_X1 \EXU/CSRControl/_2600_ ( .A(\EXU/CSRControl/_0624_ ), .B1(\EXU/CSRControl/_0369_ ), .B2(\EXU/CSRControl/_0625_ ), .ZN(\EXU/CSRControl/_0654_ ) );
AOI21_X1 \EXU/CSRControl/_2601_ ( .A(\EXU/CSRControl/_0652_ ), .B1(\EXU/CSRControl/_0653_ ), .B2(\EXU/CSRControl/_0654_ ), .ZN(\EXU/CSRControl/_0076_ ) );
OAI21_X1 \EXU/CSRControl/_2602_ ( .A(\EXU/CSRControl/_0648_ ), .B1(\EXU/CSRControl/_0619_ ), .B2(\EXU/CSRControl/_0227_ ), .ZN(\EXU/CSRControl/_0655_ ) );
AND2_X1 \EXU/CSRControl/_2603_ ( .A1(\EXU/CSRControl/_1328_ ), .A2(\EXU/CSRControl/_1329_ ), .ZN(\EXU/CSRControl/_0656_ ) );
OR2_X1 \EXU/CSRControl/_2604_ ( .A1(\EXU/CSRControl/_0656_ ), .A2(\EXU/CSRControl/_0645_ ), .ZN(\EXU/CSRControl/_0657_ ) );
AOI21_X1 \EXU/CSRControl/_2605_ ( .A(\EXU/CSRControl/_0624_ ), .B1(\EXU/CSRControl/_0370_ ), .B2(\EXU/CSRControl/_0625_ ), .ZN(\EXU/CSRControl/_0658_ ) );
AOI21_X1 \EXU/CSRControl/_2606_ ( .A(\EXU/CSRControl/_0655_ ), .B1(\EXU/CSRControl/_0657_ ), .B2(\EXU/CSRControl/_0658_ ), .ZN(\EXU/CSRControl/_0077_ ) );
BUF_X4 \EXU/CSRControl/_2607_ ( .A(\EXU/CSRControl/_0618_ ), .Z(\EXU/CSRControl/_0659_ ) );
OAI21_X1 \EXU/CSRControl/_2608_ ( .A(\EXU/CSRControl/_0648_ ), .B1(\EXU/CSRControl/_0659_ ), .B2(\EXU/CSRControl/_0197_ ), .ZN(\EXU/CSRControl/_0660_ ) );
AND2_X1 \EXU/CSRControl/_2609_ ( .A1(\EXU/CSRControl/_1339_ ), .A2(\EXU/CSRControl/_1340_ ), .ZN(\EXU/CSRControl/_0661_ ) );
OR2_X1 \EXU/CSRControl/_2610_ ( .A1(\EXU/CSRControl/_0661_ ), .A2(\EXU/CSRControl/_0645_ ), .ZN(\EXU/CSRControl/_0662_ ) );
BUF_X4 \EXU/CSRControl/_2611_ ( .A(\EXU/CSRControl/_0623_ ), .Z(\EXU/CSRControl/_0663_ ) );
BUF_X4 \EXU/CSRControl/_2612_ ( .A(\EXU/CSRControl/_1160_ ), .Z(\EXU/CSRControl/_0664_ ) );
AOI21_X1 \EXU/CSRControl/_2613_ ( .A(\EXU/CSRControl/_0663_ ), .B1(\EXU/CSRControl/_0340_ ), .B2(\EXU/CSRControl/_0664_ ), .ZN(\EXU/CSRControl/_0665_ ) );
AOI21_X1 \EXU/CSRControl/_2614_ ( .A(\EXU/CSRControl/_0660_ ), .B1(\EXU/CSRControl/_0662_ ), .B2(\EXU/CSRControl/_0665_ ), .ZN(\EXU/CSRControl/_0078_ ) );
OAI21_X1 \EXU/CSRControl/_2615_ ( .A(\EXU/CSRControl/_0648_ ), .B1(\EXU/CSRControl/_0659_ ), .B2(\EXU/CSRControl/_0198_ ), .ZN(\EXU/CSRControl/_0666_ ) );
INV_X1 \EXU/CSRControl/_2616_ ( .A(\EXU/CSRControl/_1199_ ), .ZN(\EXU/CSRControl/_0667_ ) );
AOI21_X1 \EXU/CSRControl/_2617_ ( .A(\EXU/CSRControl/_0663_ ), .B1(\EXU/CSRControl/_0341_ ), .B2(\EXU/CSRControl/_0664_ ), .ZN(\EXU/CSRControl/_0668_ ) );
AOI21_X1 \EXU/CSRControl/_2618_ ( .A(\EXU/CSRControl/_0666_ ), .B1(\EXU/CSRControl/_0667_ ), .B2(\EXU/CSRControl/_0668_ ), .ZN(\EXU/CSRControl/_0079_ ) );
OAI21_X1 \EXU/CSRControl/_2619_ ( .A(\EXU/CSRControl/_0648_ ), .B1(\EXU/CSRControl/_0659_ ), .B2(\EXU/CSRControl/_0199_ ), .ZN(\EXU/CSRControl/_0669_ ) );
AND2_X2 \EXU/CSRControl/_2620_ ( .A1(\EXU/CSRControl/_1216_ ), .A2(\EXU/CSRControl/_1217_ ), .ZN(\EXU/CSRControl/_0670_ ) );
OR2_X4 \EXU/CSRControl/_2621_ ( .A1(\EXU/CSRControl/_0670_ ), .A2(\EXU/CSRControl/_0645_ ), .ZN(\EXU/CSRControl/_0671_ ) );
AOI21_X1 \EXU/CSRControl/_2622_ ( .A(\EXU/CSRControl/_0663_ ), .B1(\EXU/CSRControl/_0342_ ), .B2(\EXU/CSRControl/_0664_ ), .ZN(\EXU/CSRControl/_0672_ ) );
AOI21_X1 \EXU/CSRControl/_2623_ ( .A(\EXU/CSRControl/_0669_ ), .B1(\EXU/CSRControl/_0671_ ), .B2(\EXU/CSRControl/_0672_ ), .ZN(\EXU/CSRControl/_0080_ ) );
OAI21_X1 \EXU/CSRControl/_2624_ ( .A(\EXU/CSRControl/_0648_ ), .B1(\EXU/CSRControl/_0659_ ), .B2(\EXU/CSRControl/_0200_ ), .ZN(\EXU/CSRControl/_0673_ ) );
AND2_X1 \EXU/CSRControl/_2625_ ( .A1(\EXU/CSRControl/_1349_ ), .A2(\EXU/CSRControl/_1350_ ), .ZN(\EXU/CSRControl/_0674_ ) );
OR2_X2 \EXU/CSRControl/_2626_ ( .A1(\EXU/CSRControl/_0674_ ), .A2(\EXU/CSRControl/_0645_ ), .ZN(\EXU/CSRControl/_0675_ ) );
AOI21_X1 \EXU/CSRControl/_2627_ ( .A(\EXU/CSRControl/_0663_ ), .B1(\EXU/CSRControl/_0343_ ), .B2(\EXU/CSRControl/_0664_ ), .ZN(\EXU/CSRControl/_0676_ ) );
AOI21_X1 \EXU/CSRControl/_2628_ ( .A(\EXU/CSRControl/_0673_ ), .B1(\EXU/CSRControl/_0675_ ), .B2(\EXU/CSRControl/_0676_ ), .ZN(\EXU/CSRControl/_0081_ ) );
OAI21_X1 \EXU/CSRControl/_2629_ ( .A(\EXU/CSRControl/_0648_ ), .B1(\EXU/CSRControl/_0659_ ), .B2(\EXU/CSRControl/_0201_ ), .ZN(\EXU/CSRControl/_0677_ ) );
OR2_X1 \EXU/CSRControl/_2630_ ( .A1(\EXU/CSRControl/_1361_ ), .A2(\EXU/CSRControl/_0645_ ), .ZN(\EXU/CSRControl/_0678_ ) );
AOI21_X1 \EXU/CSRControl/_2631_ ( .A(\EXU/CSRControl/_0663_ ), .B1(\EXU/CSRControl/_0344_ ), .B2(\EXU/CSRControl/_0664_ ), .ZN(\EXU/CSRControl/_0679_ ) );
AOI21_X1 \EXU/CSRControl/_2632_ ( .A(\EXU/CSRControl/_0677_ ), .B1(\EXU/CSRControl/_0678_ ), .B2(\EXU/CSRControl/_0679_ ), .ZN(\EXU/CSRControl/_0082_ ) );
OAI21_X1 \EXU/CSRControl/_2633_ ( .A(\EXU/CSRControl/_0648_ ), .B1(\EXU/CSRControl/_0659_ ), .B2(\EXU/CSRControl/_0202_ ), .ZN(\EXU/CSRControl/_0680_ ) );
AND2_X1 \EXU/CSRControl/_2634_ ( .A1(\EXU/CSRControl/_1369_ ), .A2(\EXU/CSRControl/_1370_ ), .ZN(\EXU/CSRControl/_0681_ ) );
OR2_X4 \EXU/CSRControl/_2635_ ( .A1(\EXU/CSRControl/_0681_ ), .A2(\EXU/CSRControl/_0645_ ), .ZN(\EXU/CSRControl/_0682_ ) );
AOI21_X1 \EXU/CSRControl/_2636_ ( .A(\EXU/CSRControl/_0663_ ), .B1(\EXU/CSRControl/_0345_ ), .B2(\EXU/CSRControl/_0664_ ), .ZN(\EXU/CSRControl/_0683_ ) );
AOI21_X1 \EXU/CSRControl/_2637_ ( .A(\EXU/CSRControl/_0680_ ), .B1(\EXU/CSRControl/_0682_ ), .B2(\EXU/CSRControl/_0683_ ), .ZN(\EXU/CSRControl/_0083_ ) );
OAI21_X1 \EXU/CSRControl/_2638_ ( .A(\EXU/CSRControl/_0648_ ), .B1(\EXU/CSRControl/_0659_ ), .B2(\EXU/CSRControl/_0203_ ), .ZN(\EXU/CSRControl/_0684_ ) );
OR2_X2 \EXU/CSRControl/_2639_ ( .A1(\EXU/CSRControl/_0382_ ), .A2(\EXU/CSRControl/_0645_ ), .ZN(\EXU/CSRControl/_0685_ ) );
AOI21_X1 \EXU/CSRControl/_2640_ ( .A(\EXU/CSRControl/_0663_ ), .B1(\EXU/CSRControl/_0346_ ), .B2(\EXU/CSRControl/_0664_ ), .ZN(\EXU/CSRControl/_0686_ ) );
AOI21_X1 \EXU/CSRControl/_2641_ ( .A(\EXU/CSRControl/_0684_ ), .B1(\EXU/CSRControl/_0685_ ), .B2(\EXU/CSRControl/_0686_ ), .ZN(\EXU/CSRControl/_0084_ ) );
BUF_X4 \EXU/CSRControl/_2642_ ( .A(\EXU/CSRControl/_1221_ ), .Z(\EXU/CSRControl/_0687_ ) );
OAI21_X1 \EXU/CSRControl/_2643_ ( .A(\EXU/CSRControl/_0687_ ), .B1(\EXU/CSRControl/_0659_ ), .B2(\EXU/CSRControl/_0204_ ), .ZN(\EXU/CSRControl/_0688_ ) );
AND2_X1 \EXU/CSRControl/_2644_ ( .A1(\EXU/CSRControl/_0391_ ), .A2(\EXU/CSRControl/_0392_ ), .ZN(\EXU/CSRControl/_0689_ ) );
CLKBUF_X2 \EXU/CSRControl/_2645_ ( .A(\EXU/CSRControl/_0841_ ), .Z(\EXU/CSRControl/_0690_ ) );
OR2_X1 \EXU/CSRControl/_2646_ ( .A1(\EXU/CSRControl/_0689_ ), .A2(\EXU/CSRControl/_0690_ ), .ZN(\EXU/CSRControl/_0691_ ) );
AOI21_X1 \EXU/CSRControl/_2647_ ( .A(\EXU/CSRControl/_0663_ ), .B1(\EXU/CSRControl/_0347_ ), .B2(\EXU/CSRControl/_0664_ ), .ZN(\EXU/CSRControl/_0692_ ) );
AOI21_X1 \EXU/CSRControl/_2648_ ( .A(\EXU/CSRControl/_0688_ ), .B1(\EXU/CSRControl/_0691_ ), .B2(\EXU/CSRControl/_0692_ ), .ZN(\EXU/CSRControl/_0085_ ) );
OAI21_X1 \EXU/CSRControl/_2649_ ( .A(\EXU/CSRControl/_0687_ ), .B1(\EXU/CSRControl/_0659_ ), .B2(\EXU/CSRControl/_0205_ ), .ZN(\EXU/CSRControl/_0693_ ) );
AND2_X1 \EXU/CSRControl/_2650_ ( .A1(\EXU/CSRControl/_0402_ ), .A2(\EXU/CSRControl/_0403_ ), .ZN(\EXU/CSRControl/_0694_ ) );
OR2_X1 \EXU/CSRControl/_2651_ ( .A1(\EXU/CSRControl/_0694_ ), .A2(\EXU/CSRControl/_0690_ ), .ZN(\EXU/CSRControl/_0695_ ) );
AOI21_X1 \EXU/CSRControl/_2652_ ( .A(\EXU/CSRControl/_0663_ ), .B1(\EXU/CSRControl/_0348_ ), .B2(\EXU/CSRControl/_0664_ ), .ZN(\EXU/CSRControl/_0696_ ) );
AOI21_X1 \EXU/CSRControl/_2653_ ( .A(\EXU/CSRControl/_0693_ ), .B1(\EXU/CSRControl/_0695_ ), .B2(\EXU/CSRControl/_0696_ ), .ZN(\EXU/CSRControl/_0086_ ) );
OAI21_X1 \EXU/CSRControl/_2654_ ( .A(\EXU/CSRControl/_0687_ ), .B1(\EXU/CSRControl/_0659_ ), .B2(\EXU/CSRControl/_0206_ ), .ZN(\EXU/CSRControl/_0697_ ) );
OR2_X2 \EXU/CSRControl/_2655_ ( .A1(\EXU/CSRControl/_0415_ ), .A2(\EXU/CSRControl/_0690_ ), .ZN(\EXU/CSRControl/_0698_ ) );
AOI21_X1 \EXU/CSRControl/_2656_ ( .A(\EXU/CSRControl/_0663_ ), .B1(\EXU/CSRControl/_0349_ ), .B2(\EXU/CSRControl/_0664_ ), .ZN(\EXU/CSRControl/_0699_ ) );
AOI21_X1 \EXU/CSRControl/_2657_ ( .A(\EXU/CSRControl/_0697_ ), .B1(\EXU/CSRControl/_0698_ ), .B2(\EXU/CSRControl/_0699_ ), .ZN(\EXU/CSRControl/_0087_ ) );
BUF_X4 \EXU/CSRControl/_2658_ ( .A(\EXU/CSRControl/_0618_ ), .Z(\EXU/CSRControl/_0700_ ) );
OAI21_X1 \EXU/CSRControl/_2659_ ( .A(\EXU/CSRControl/_0687_ ), .B1(\EXU/CSRControl/_0700_ ), .B2(\EXU/CSRControl/_0208_ ), .ZN(\EXU/CSRControl/_0701_ ) );
OR2_X2 \EXU/CSRControl/_2660_ ( .A1(\EXU/CSRControl/_0426_ ), .A2(\EXU/CSRControl/_0690_ ), .ZN(\EXU/CSRControl/_0702_ ) );
BUF_X4 \EXU/CSRControl/_2661_ ( .A(\EXU/CSRControl/_0623_ ), .Z(\EXU/CSRControl/_0703_ ) );
BUF_X4 \EXU/CSRControl/_2662_ ( .A(\EXU/CSRControl/_0841_ ), .Z(\EXU/CSRControl/_0704_ ) );
AOI21_X1 \EXU/CSRControl/_2663_ ( .A(\EXU/CSRControl/_0703_ ), .B1(\EXU/CSRControl/_0351_ ), .B2(\EXU/CSRControl/_0704_ ), .ZN(\EXU/CSRControl/_0705_ ) );
AOI21_X1 \EXU/CSRControl/_2664_ ( .A(\EXU/CSRControl/_0701_ ), .B1(\EXU/CSRControl/_0702_ ), .B2(\EXU/CSRControl/_0705_ ), .ZN(\EXU/CSRControl/_0088_ ) );
OAI21_X1 \EXU/CSRControl/_2665_ ( .A(\EXU/CSRControl/_0687_ ), .B1(\EXU/CSRControl/_0700_ ), .B2(\EXU/CSRControl/_0209_ ), .ZN(\EXU/CSRControl/_0706_ ) );
OR2_X4 \EXU/CSRControl/_2666_ ( .A1(\EXU/CSRControl/_0436_ ), .A2(\EXU/CSRControl/_0690_ ), .ZN(\EXU/CSRControl/_0707_ ) );
AOI21_X1 \EXU/CSRControl/_2667_ ( .A(\EXU/CSRControl/_0703_ ), .B1(\EXU/CSRControl/_0352_ ), .B2(\EXU/CSRControl/_0704_ ), .ZN(\EXU/CSRControl/_0708_ ) );
AOI21_X1 \EXU/CSRControl/_2668_ ( .A(\EXU/CSRControl/_0706_ ), .B1(\EXU/CSRControl/_0707_ ), .B2(\EXU/CSRControl/_0708_ ), .ZN(\EXU/CSRControl/_0089_ ) );
OAI21_X1 \EXU/CSRControl/_2669_ ( .A(\EXU/CSRControl/_0687_ ), .B1(\EXU/CSRControl/_0700_ ), .B2(\EXU/CSRControl/_0210_ ), .ZN(\EXU/CSRControl/_0709_ ) );
AND2_X1 \EXU/CSRControl/_2670_ ( .A1(\EXU/CSRControl/_0442_ ), .A2(\EXU/CSRControl/_0443_ ), .ZN(\EXU/CSRControl/_0710_ ) );
OR2_X1 \EXU/CSRControl/_2671_ ( .A1(\EXU/CSRControl/_0710_ ), .A2(\EXU/CSRControl/_0690_ ), .ZN(\EXU/CSRControl/_0711_ ) );
AOI21_X1 \EXU/CSRControl/_2672_ ( .A(\EXU/CSRControl/_0703_ ), .B1(\EXU/CSRControl/_0353_ ), .B2(\EXU/CSRControl/_0704_ ), .ZN(\EXU/CSRControl/_0712_ ) );
AOI21_X1 \EXU/CSRControl/_2673_ ( .A(\EXU/CSRControl/_0709_ ), .B1(\EXU/CSRControl/_0711_ ), .B2(\EXU/CSRControl/_0712_ ), .ZN(\EXU/CSRControl/_0090_ ) );
OAI21_X1 \EXU/CSRControl/_2674_ ( .A(\EXU/CSRControl/_0687_ ), .B1(\EXU/CSRControl/_0700_ ), .B2(\EXU/CSRControl/_0211_ ), .ZN(\EXU/CSRControl/_0713_ ) );
AND2_X1 \EXU/CSRControl/_2675_ ( .A1(\EXU/CSRControl/_0453_ ), .A2(\EXU/CSRControl/_0454_ ), .ZN(\EXU/CSRControl/_0714_ ) );
OR2_X1 \EXU/CSRControl/_2676_ ( .A1(\EXU/CSRControl/_0714_ ), .A2(\EXU/CSRControl/_0690_ ), .ZN(\EXU/CSRControl/_0715_ ) );
AOI21_X1 \EXU/CSRControl/_2677_ ( .A(\EXU/CSRControl/_0703_ ), .B1(\EXU/CSRControl/_0354_ ), .B2(\EXU/CSRControl/_0704_ ), .ZN(\EXU/CSRControl/_0716_ ) );
AOI21_X1 \EXU/CSRControl/_2678_ ( .A(\EXU/CSRControl/_0713_ ), .B1(\EXU/CSRControl/_0715_ ), .B2(\EXU/CSRControl/_0716_ ), .ZN(\EXU/CSRControl/_0091_ ) );
OAI21_X1 \EXU/CSRControl/_2679_ ( .A(\EXU/CSRControl/_0687_ ), .B1(\EXU/CSRControl/_0700_ ), .B2(\EXU/CSRControl/_0212_ ), .ZN(\EXU/CSRControl/_0717_ ) );
OR2_X4 \EXU/CSRControl/_2680_ ( .A1(\EXU/CSRControl/_0467_ ), .A2(\EXU/CSRControl/_0690_ ), .ZN(\EXU/CSRControl/_0718_ ) );
AOI21_X1 \EXU/CSRControl/_2681_ ( .A(\EXU/CSRControl/_0703_ ), .B1(\EXU/CSRControl/_0355_ ), .B2(\EXU/CSRControl/_0704_ ), .ZN(\EXU/CSRControl/_0719_ ) );
AOI21_X1 \EXU/CSRControl/_2682_ ( .A(\EXU/CSRControl/_0717_ ), .B1(\EXU/CSRControl/_0718_ ), .B2(\EXU/CSRControl/_0719_ ), .ZN(\EXU/CSRControl/_0092_ ) );
OAI21_X1 \EXU/CSRControl/_2683_ ( .A(\EXU/CSRControl/_0687_ ), .B1(\EXU/CSRControl/_0700_ ), .B2(\EXU/CSRControl/_0213_ ), .ZN(\EXU/CSRControl/_0720_ ) );
AND2_X1 \EXU/CSRControl/_2684_ ( .A1(\EXU/CSRControl/_0475_ ), .A2(\EXU/CSRControl/_0476_ ), .ZN(\EXU/CSRControl/_0721_ ) );
OR2_X1 \EXU/CSRControl/_2685_ ( .A1(\EXU/CSRControl/_0721_ ), .A2(\EXU/CSRControl/_0690_ ), .ZN(\EXU/CSRControl/_0722_ ) );
AOI21_X1 \EXU/CSRControl/_2686_ ( .A(\EXU/CSRControl/_0703_ ), .B1(\EXU/CSRControl/_0356_ ), .B2(\EXU/CSRControl/_0704_ ), .ZN(\EXU/CSRControl/_0723_ ) );
AOI21_X1 \EXU/CSRControl/_2687_ ( .A(\EXU/CSRControl/_0720_ ), .B1(\EXU/CSRControl/_0722_ ), .B2(\EXU/CSRControl/_0723_ ), .ZN(\EXU/CSRControl/_0093_ ) );
OAI21_X1 \EXU/CSRControl/_2688_ ( .A(\EXU/CSRControl/_0687_ ), .B1(\EXU/CSRControl/_0700_ ), .B2(\EXU/CSRControl/_0214_ ), .ZN(\EXU/CSRControl/_0724_ ) );
AND2_X1 \EXU/CSRControl/_2689_ ( .A1(\EXU/CSRControl/_0487_ ), .A2(\EXU/CSRControl/_0488_ ), .ZN(\EXU/CSRControl/_0725_ ) );
OR2_X1 \EXU/CSRControl/_2690_ ( .A1(\EXU/CSRControl/_0725_ ), .A2(\EXU/CSRControl/_0690_ ), .ZN(\EXU/CSRControl/_0726_ ) );
AOI21_X1 \EXU/CSRControl/_2691_ ( .A(\EXU/CSRControl/_0703_ ), .B1(\EXU/CSRControl/_0357_ ), .B2(\EXU/CSRControl/_0704_ ), .ZN(\EXU/CSRControl/_0727_ ) );
AOI21_X1 \EXU/CSRControl/_2692_ ( .A(\EXU/CSRControl/_0724_ ), .B1(\EXU/CSRControl/_0726_ ), .B2(\EXU/CSRControl/_0727_ ), .ZN(\EXU/CSRControl/_0094_ ) );
BUF_X4 \EXU/CSRControl/_2693_ ( .A(\EXU/CSRControl/_1221_ ), .Z(\EXU/CSRControl/_0728_ ) );
OAI21_X1 \EXU/CSRControl/_2694_ ( .A(\EXU/CSRControl/_0728_ ), .B1(\EXU/CSRControl/_0700_ ), .B2(\EXU/CSRControl/_0215_ ), .ZN(\EXU/CSRControl/_0729_ ) );
AND2_X1 \EXU/CSRControl/_2695_ ( .A1(\EXU/CSRControl/_0497_ ), .A2(\EXU/CSRControl/_0498_ ), .ZN(\EXU/CSRControl/_0730_ ) );
OR2_X2 \EXU/CSRControl/_2696_ ( .A1(\EXU/CSRControl/_0730_ ), .A2(\EXU/CSRControl/_1160_ ), .ZN(\EXU/CSRControl/_0731_ ) );
AOI21_X1 \EXU/CSRControl/_2697_ ( .A(\EXU/CSRControl/_0703_ ), .B1(\EXU/CSRControl/_0358_ ), .B2(\EXU/CSRControl/_0704_ ), .ZN(\EXU/CSRControl/_0732_ ) );
AOI21_X1 \EXU/CSRControl/_2698_ ( .A(\EXU/CSRControl/_0729_ ), .B1(\EXU/CSRControl/_0731_ ), .B2(\EXU/CSRControl/_0732_ ), .ZN(\EXU/CSRControl/_0095_ ) );
OAI21_X1 \EXU/CSRControl/_2699_ ( .A(\EXU/CSRControl/_0728_ ), .B1(\EXU/CSRControl/_0700_ ), .B2(\EXU/CSRControl/_0216_ ), .ZN(\EXU/CSRControl/_0733_ ) );
AND2_X1 \EXU/CSRControl/_2700_ ( .A1(\EXU/CSRControl/_0507_ ), .A2(\EXU/CSRControl/_0508_ ), .ZN(\EXU/CSRControl/_0734_ ) );
OR2_X1 \EXU/CSRControl/_2701_ ( .A1(\EXU/CSRControl/_0734_ ), .A2(\EXU/CSRControl/_1160_ ), .ZN(\EXU/CSRControl/_0735_ ) );
AOI21_X1 \EXU/CSRControl/_2702_ ( .A(\EXU/CSRControl/_0703_ ), .B1(\EXU/CSRControl/_0359_ ), .B2(\EXU/CSRControl/_0704_ ), .ZN(\EXU/CSRControl/_0736_ ) );
AOI21_X1 \EXU/CSRControl/_2703_ ( .A(\EXU/CSRControl/_0733_ ), .B1(\EXU/CSRControl/_0735_ ), .B2(\EXU/CSRControl/_0736_ ), .ZN(\EXU/CSRControl/_0096_ ) );
OAI21_X1 \EXU/CSRControl/_2704_ ( .A(\EXU/CSRControl/_0728_ ), .B1(\EXU/CSRControl/_0700_ ), .B2(\EXU/CSRControl/_0217_ ), .ZN(\EXU/CSRControl/_0737_ ) );
OR2_X2 \EXU/CSRControl/_2705_ ( .A1(\EXU/CSRControl/_0520_ ), .A2(\EXU/CSRControl/_1160_ ), .ZN(\EXU/CSRControl/_0738_ ) );
AOI21_X1 \EXU/CSRControl/_2706_ ( .A(\EXU/CSRControl/_0703_ ), .B1(\EXU/CSRControl/_0360_ ), .B2(\EXU/CSRControl/_0704_ ), .ZN(\EXU/CSRControl/_0739_ ) );
AOI21_X1 \EXU/CSRControl/_2707_ ( .A(\EXU/CSRControl/_0737_ ), .B1(\EXU/CSRControl/_0738_ ), .B2(\EXU/CSRControl/_0739_ ), .ZN(\EXU/CSRControl/_0097_ ) );
OAI21_X1 \EXU/CSRControl/_2708_ ( .A(\EXU/CSRControl/_0728_ ), .B1(\EXU/CSRControl/_0618_ ), .B2(\EXU/CSRControl/_0219_ ), .ZN(\EXU/CSRControl/_0740_ ) );
OR2_X1 \EXU/CSRControl/_2709_ ( .A1(\EXU/CSRControl/_0530_ ), .A2(\EXU/CSRControl/_1160_ ), .ZN(\EXU/CSRControl/_0741_ ) );
AOI21_X1 \EXU/CSRControl/_2710_ ( .A(\EXU/CSRControl/_0623_ ), .B1(\EXU/CSRControl/_0362_ ), .B2(\EXU/CSRControl/_1200_ ), .ZN(\EXU/CSRControl/_0742_ ) );
AOI21_X1 \EXU/CSRControl/_2711_ ( .A(\EXU/CSRControl/_0740_ ), .B1(\EXU/CSRControl/_0741_ ), .B2(\EXU/CSRControl/_0742_ ), .ZN(\EXU/CSRControl/_0098_ ) );
OAI21_X1 \EXU/CSRControl/_2712_ ( .A(\EXU/CSRControl/_0728_ ), .B1(\EXU/CSRControl/_0618_ ), .B2(\EXU/CSRControl/_0220_ ), .ZN(\EXU/CSRControl/_0743_ ) );
AND2_X1 \EXU/CSRControl/_2713_ ( .A1(\EXU/CSRControl/_0539_ ), .A2(\EXU/CSRControl/_0540_ ), .ZN(\EXU/CSRControl/_0744_ ) );
OR2_X1 \EXU/CSRControl/_2714_ ( .A1(\EXU/CSRControl/_0744_ ), .A2(\EXU/CSRControl/_1160_ ), .ZN(\EXU/CSRControl/_0745_ ) );
AOI21_X1 \EXU/CSRControl/_2715_ ( .A(\EXU/CSRControl/_0623_ ), .B1(\EXU/CSRControl/_0363_ ), .B2(\EXU/CSRControl/_1200_ ), .ZN(\EXU/CSRControl/_0746_ ) );
AOI21_X1 \EXU/CSRControl/_2716_ ( .A(\EXU/CSRControl/_0743_ ), .B1(\EXU/CSRControl/_0745_ ), .B2(\EXU/CSRControl/_0746_ ), .ZN(\EXU/CSRControl/_0099_ ) );
OR2_X4 \EXU/CSRControl/_2717_ ( .A1(\EXU/CSRControl/_1205_ ), .A2(\EXU/CSRControl/_0795_ ), .ZN(\EXU/CSRControl/_0747_ ) );
AND2_X2 \EXU/CSRControl/_2718_ ( .A1(\EXU/CSRControl/_0747_ ), .A2(\EXU/CSRControl/_0617_ ), .ZN(\EXU/CSRControl/_0748_ ) );
BUF_X8 \EXU/CSRControl/_2719_ ( .A(\EXU/CSRControl/_0748_ ), .Z(\EXU/CSRControl/_0749_ ) );
BUF_X4 \EXU/CSRControl/_2720_ ( .A(\EXU/CSRControl/_0749_ ), .Z(\EXU/CSRControl/_0750_ ) );
OAI21_X1 \EXU/CSRControl/_2721_ ( .A(\EXU/CSRControl/_0728_ ), .B1(\EXU/CSRControl/_0750_ ), .B2(\EXU/CSRControl/_0132_ ), .ZN(\EXU/CSRControl/_0751_ ) );
INV_X4 \EXU/CSRControl/_2722_ ( .A(\EXU/CSRControl/_0749_ ), .ZN(\EXU/CSRControl/_0752_ ) );
AOI21_X1 \EXU/CSRControl/_2723_ ( .A(\EXU/CSRControl/_0752_ ), .B1(\EXU/CSRControl/_1372_ ), .B2(\EXU/CSRControl/_1200_ ), .ZN(\EXU/CSRControl/_0753_ ) );
AOI21_X1 \EXU/CSRControl/_2724_ ( .A(\EXU/CSRControl/_0751_ ), .B1(\EXU/CSRControl/_0622_ ), .B2(\EXU/CSRControl/_0753_ ), .ZN(\EXU/CSRControl/_0100_ ) );
BUF_X4 \EXU/CSRControl/_2725_ ( .A(\EXU/CSRControl/_0749_ ), .Z(\EXU/CSRControl/_0754_ ) );
OAI21_X1 \EXU/CSRControl/_2726_ ( .A(\EXU/CSRControl/_0728_ ), .B1(\EXU/CSRControl/_0754_ ), .B2(\EXU/CSRControl/_0143_ ), .ZN(\EXU/CSRControl/_0755_ ) );
NOR2_X1 \EXU/CSRControl/_2727_ ( .A1(\EXU/CSRControl/_0752_ ), .A2(\EXU/CSRControl/_1219_ ), .ZN(\EXU/CSRControl/_0756_ ) );
AOI21_X1 \EXU/CSRControl/_2728_ ( .A(\EXU/CSRControl/_0755_ ), .B1(\EXU/CSRControl/_0629_ ), .B2(\EXU/CSRControl/_0756_ ), .ZN(\EXU/CSRControl/_0101_ ) );
OAI21_X1 \EXU/CSRControl/_2729_ ( .A(\EXU/CSRControl/_0728_ ), .B1(\EXU/CSRControl/_0754_ ), .B2(\EXU/CSRControl/_0154_ ), .ZN(\EXU/CSRControl/_0757_ ) );
BUF_X4 \EXU/CSRControl/_2730_ ( .A(\EXU/CSRControl/_0749_ ), .Z(\EXU/CSRControl/_0758_ ) );
AOI21_X1 \EXU/CSRControl/_2731_ ( .A(\EXU/CSRControl/_0757_ ), .B1(\EXU/CSRControl/_0632_ ), .B2(\EXU/CSRControl/_0758_ ), .ZN(\EXU/CSRControl/_0102_ ) );
OAI21_X1 \EXU/CSRControl/_2732_ ( .A(\EXU/CSRControl/_0728_ ), .B1(\EXU/CSRControl/_0754_ ), .B2(\EXU/CSRControl/_0157_ ), .ZN(\EXU/CSRControl/_0759_ ) );
NOR4_X1 \EXU/CSRControl/_2733_ ( .A1(\EXU/CSRControl/_0800_ ), .A2(\EXU/CSRControl/_0273_ ), .A3(\EXU/CSRControl/_0272_ ), .A4(\EXU/CSRControl/_1373_ ), .ZN(\EXU/CSRControl/_0760_ ) );
AOI211_X2 \EXU/CSRControl/_2734_ ( .A(\EXU/CSRControl/_0760_ ), .B(\EXU/CSRControl/_0752_ ), .C1(\EXU/CSRControl/_1372_ ), .C2(\EXU/CSRControl/_0841_ ), .ZN(\EXU/CSRControl/_0761_ ) );
AOI21_X1 \EXU/CSRControl/_2735_ ( .A(\EXU/CSRControl/_0759_ ), .B1(\EXU/CSRControl/_0761_ ), .B2(\EXU/CSRControl/_0635_ ), .ZN(\EXU/CSRControl/_0103_ ) );
OAI21_X1 \EXU/CSRControl/_2736_ ( .A(\EXU/CSRControl/_0728_ ), .B1(\EXU/CSRControl/_0754_ ), .B2(\EXU/CSRControl/_0158_ ), .ZN(\EXU/CSRControl/_0762_ ) );
AOI21_X1 \EXU/CSRControl/_2737_ ( .A(\EXU/CSRControl/_0762_ ), .B1(\EXU/CSRControl/_0638_ ), .B2(\EXU/CSRControl/_0758_ ), .ZN(\EXU/CSRControl/_0104_ ) );
BUF_X4 \EXU/CSRControl/_2738_ ( .A(\EXU/CSRControl/_1221_ ), .Z(\EXU/CSRControl/_0763_ ) );
OAI21_X1 \EXU/CSRControl/_2739_ ( .A(\EXU/CSRControl/_0763_ ), .B1(\EXU/CSRControl/_0754_ ), .B2(\EXU/CSRControl/_0159_ ), .ZN(\EXU/CSRControl/_0764_ ) );
AOI21_X1 \EXU/CSRControl/_2740_ ( .A(\EXU/CSRControl/_0764_ ), .B1(\EXU/CSRControl/_0641_ ), .B2(\EXU/CSRControl/_0758_ ), .ZN(\EXU/CSRControl/_0105_ ) );
OAI21_X1 \EXU/CSRControl/_2741_ ( .A(\EXU/CSRControl/_0763_ ), .B1(\EXU/CSRControl/_0754_ ), .B2(\EXU/CSRControl/_0160_ ), .ZN(\EXU/CSRControl/_0765_ ) );
AOI21_X1 \EXU/CSRControl/_2742_ ( .A(\EXU/CSRControl/_0765_ ), .B1(\EXU/CSRControl/_0646_ ), .B2(\EXU/CSRControl/_0758_ ), .ZN(\EXU/CSRControl/_0106_ ) );
OAI21_X1 \EXU/CSRControl/_2743_ ( .A(\EXU/CSRControl/_0763_ ), .B1(\EXU/CSRControl/_0754_ ), .B2(\EXU/CSRControl/_0161_ ), .ZN(\EXU/CSRControl/_0766_ ) );
AOI21_X1 \EXU/CSRControl/_2744_ ( .A(\EXU/CSRControl/_0766_ ), .B1(\EXU/CSRControl/_0650_ ), .B2(\EXU/CSRControl/_0758_ ), .ZN(\EXU/CSRControl/_0107_ ) );
OAI21_X1 \EXU/CSRControl/_2745_ ( .A(\EXU/CSRControl/_0763_ ), .B1(\EXU/CSRControl/_0754_ ), .B2(\EXU/CSRControl/_0162_ ), .ZN(\EXU/CSRControl/_0767_ ) );
AOI21_X1 \EXU/CSRControl/_2746_ ( .A(\EXU/CSRControl/_0767_ ), .B1(\EXU/CSRControl/_0653_ ), .B2(\EXU/CSRControl/_0758_ ), .ZN(\EXU/CSRControl/_0108_ ) );
OAI21_X1 \EXU/CSRControl/_2747_ ( .A(\EXU/CSRControl/_0763_ ), .B1(\EXU/CSRControl/_0754_ ), .B2(\EXU/CSRControl/_0163_ ), .ZN(\EXU/CSRControl/_0768_ ) );
AOI21_X1 \EXU/CSRControl/_2748_ ( .A(\EXU/CSRControl/_0768_ ), .B1(\EXU/CSRControl/_0657_ ), .B2(\EXU/CSRControl/_0758_ ), .ZN(\EXU/CSRControl/_0109_ ) );
OAI21_X1 \EXU/CSRControl/_2749_ ( .A(\EXU/CSRControl/_0763_ ), .B1(\EXU/CSRControl/_0754_ ), .B2(\EXU/CSRControl/_0133_ ), .ZN(\EXU/CSRControl/_0769_ ) );
AOI21_X1 \EXU/CSRControl/_2750_ ( .A(\EXU/CSRControl/_0769_ ), .B1(\EXU/CSRControl/_0662_ ), .B2(\EXU/CSRControl/_0758_ ), .ZN(\EXU/CSRControl/_0110_ ) );
BUF_X4 \EXU/CSRControl/_2751_ ( .A(\EXU/CSRControl/_0749_ ), .Z(\EXU/CSRControl/_0770_ ) );
OAI21_X1 \EXU/CSRControl/_2752_ ( .A(\EXU/CSRControl/_0763_ ), .B1(\EXU/CSRControl/_0770_ ), .B2(\EXU/CSRControl/_0134_ ), .ZN(\EXU/CSRControl/_0771_ ) );
AOI21_X1 \EXU/CSRControl/_2753_ ( .A(\EXU/CSRControl/_0771_ ), .B1(\EXU/CSRControl/_0667_ ), .B2(\EXU/CSRControl/_0758_ ), .ZN(\EXU/CSRControl/_0111_ ) );
OAI21_X1 \EXU/CSRControl/_2754_ ( .A(\EXU/CSRControl/_0763_ ), .B1(\EXU/CSRControl/_0770_ ), .B2(\EXU/CSRControl/_0135_ ), .ZN(\EXU/CSRControl/_0772_ ) );
AOI21_X1 \EXU/CSRControl/_2755_ ( .A(\EXU/CSRControl/_0772_ ), .B1(\EXU/CSRControl/_0671_ ), .B2(\EXU/CSRControl/_0758_ ), .ZN(\EXU/CSRControl/_0112_ ) );
OAI21_X1 \EXU/CSRControl/_2756_ ( .A(\EXU/CSRControl/_0763_ ), .B1(\EXU/CSRControl/_0770_ ), .B2(\EXU/CSRControl/_0136_ ), .ZN(\EXU/CSRControl/_0773_ ) );
BUF_X4 \EXU/CSRControl/_2757_ ( .A(\EXU/CSRControl/_0749_ ), .Z(\EXU/CSRControl/_0774_ ) );
AOI21_X1 \EXU/CSRControl/_2758_ ( .A(\EXU/CSRControl/_0773_ ), .B1(\EXU/CSRControl/_0675_ ), .B2(\EXU/CSRControl/_0774_ ), .ZN(\EXU/CSRControl/_0113_ ) );
OAI21_X1 \EXU/CSRControl/_2759_ ( .A(\EXU/CSRControl/_0763_ ), .B1(\EXU/CSRControl/_0770_ ), .B2(\EXU/CSRControl/_0137_ ), .ZN(\EXU/CSRControl/_0775_ ) );
AOI21_X1 \EXU/CSRControl/_2760_ ( .A(\EXU/CSRControl/_0775_ ), .B1(\EXU/CSRControl/_0678_ ), .B2(\EXU/CSRControl/_0774_ ), .ZN(\EXU/CSRControl/_0114_ ) );
BUF_X4 \EXU/CSRControl/_2761_ ( .A(\EXU/CSRControl/_1221_ ), .Z(\EXU/CSRControl/_0776_ ) );
OAI21_X1 \EXU/CSRControl/_2762_ ( .A(\EXU/CSRControl/_0776_ ), .B1(\EXU/CSRControl/_0770_ ), .B2(\EXU/CSRControl/_0138_ ), .ZN(\EXU/CSRControl/_0777_ ) );
AOI21_X1 \EXU/CSRControl/_2763_ ( .A(\EXU/CSRControl/_0777_ ), .B1(\EXU/CSRControl/_0682_ ), .B2(\EXU/CSRControl/_0774_ ), .ZN(\EXU/CSRControl/_0115_ ) );
OAI21_X1 \EXU/CSRControl/_2764_ ( .A(\EXU/CSRControl/_0776_ ), .B1(\EXU/CSRControl/_0770_ ), .B2(\EXU/CSRControl/_0139_ ), .ZN(\EXU/CSRControl/_0778_ ) );
AOI21_X1 \EXU/CSRControl/_2765_ ( .A(\EXU/CSRControl/_0778_ ), .B1(\EXU/CSRControl/_0685_ ), .B2(\EXU/CSRControl/_0774_ ), .ZN(\EXU/CSRControl/_0116_ ) );
OAI21_X1 \EXU/CSRControl/_2766_ ( .A(\EXU/CSRControl/_0776_ ), .B1(\EXU/CSRControl/_0770_ ), .B2(\EXU/CSRControl/_0140_ ), .ZN(\EXU/CSRControl/_0779_ ) );
AOI21_X1 \EXU/CSRControl/_2767_ ( .A(\EXU/CSRControl/_0779_ ), .B1(\EXU/CSRControl/_0691_ ), .B2(\EXU/CSRControl/_0774_ ), .ZN(\EXU/CSRControl/_0117_ ) );
OAI21_X1 \EXU/CSRControl/_2768_ ( .A(\EXU/CSRControl/_0776_ ), .B1(\EXU/CSRControl/_0770_ ), .B2(\EXU/CSRControl/_0141_ ), .ZN(\EXU/CSRControl/_0780_ ) );
AOI21_X1 \EXU/CSRControl/_2769_ ( .A(\EXU/CSRControl/_0780_ ), .B1(\EXU/CSRControl/_0695_ ), .B2(\EXU/CSRControl/_0774_ ), .ZN(\EXU/CSRControl/_0118_ ) );
OAI21_X1 \EXU/CSRControl/_2770_ ( .A(\EXU/CSRControl/_0776_ ), .B1(\EXU/CSRControl/_0770_ ), .B2(\EXU/CSRControl/_0142_ ), .ZN(\EXU/CSRControl/_0781_ ) );
AOI21_X1 \EXU/CSRControl/_2771_ ( .A(\EXU/CSRControl/_0781_ ), .B1(\EXU/CSRControl/_0698_ ), .B2(\EXU/CSRControl/_0774_ ), .ZN(\EXU/CSRControl/_0119_ ) );
OAI21_X1 \EXU/CSRControl/_2772_ ( .A(\EXU/CSRControl/_0776_ ), .B1(\EXU/CSRControl/_0770_ ), .B2(\EXU/CSRControl/_0144_ ), .ZN(\EXU/CSRControl/_0782_ ) );
AOI21_X1 \EXU/CSRControl/_2773_ ( .A(\EXU/CSRControl/_0782_ ), .B1(\EXU/CSRControl/_0702_ ), .B2(\EXU/CSRControl/_0774_ ), .ZN(\EXU/CSRControl/_0120_ ) );
BUF_X4 \EXU/CSRControl/_2774_ ( .A(\EXU/CSRControl/_0749_ ), .Z(\EXU/CSRControl/_0783_ ) );
OAI21_X1 \EXU/CSRControl/_2775_ ( .A(\EXU/CSRControl/_0776_ ), .B1(\EXU/CSRControl/_0783_ ), .B2(\EXU/CSRControl/_0145_ ), .ZN(\EXU/CSRControl/_0784_ ) );
AOI21_X1 \EXU/CSRControl/_2776_ ( .A(\EXU/CSRControl/_0784_ ), .B1(\EXU/CSRControl/_0707_ ), .B2(\EXU/CSRControl/_0774_ ), .ZN(\EXU/CSRControl/_0121_ ) );
OAI21_X1 \EXU/CSRControl/_2777_ ( .A(\EXU/CSRControl/_0776_ ), .B1(\EXU/CSRControl/_0783_ ), .B2(\EXU/CSRControl/_0146_ ), .ZN(\EXU/CSRControl/_0785_ ) );
AOI21_X1 \EXU/CSRControl/_2778_ ( .A(\EXU/CSRControl/_0785_ ), .B1(\EXU/CSRControl/_0711_ ), .B2(\EXU/CSRControl/_0774_ ), .ZN(\EXU/CSRControl/_0122_ ) );
OAI21_X1 \EXU/CSRControl/_2779_ ( .A(\EXU/CSRControl/_0776_ ), .B1(\EXU/CSRControl/_0783_ ), .B2(\EXU/CSRControl/_0147_ ), .ZN(\EXU/CSRControl/_0786_ ) );
AOI21_X1 \EXU/CSRControl/_2780_ ( .A(\EXU/CSRControl/_0786_ ), .B1(\EXU/CSRControl/_0715_ ), .B2(\EXU/CSRControl/_0750_ ), .ZN(\EXU/CSRControl/_0123_ ) );
OAI21_X1 \EXU/CSRControl/_2781_ ( .A(\EXU/CSRControl/_0776_ ), .B1(\EXU/CSRControl/_0783_ ), .B2(\EXU/CSRControl/_0148_ ), .ZN(\EXU/CSRControl/_0787_ ) );
AOI21_X1 \EXU/CSRControl/_2782_ ( .A(\EXU/CSRControl/_0787_ ), .B1(\EXU/CSRControl/_0718_ ), .B2(\EXU/CSRControl/_0750_ ), .ZN(\EXU/CSRControl/_0124_ ) );
OAI21_X1 \EXU/CSRControl/_2783_ ( .A(\EXU/CSRControl/_1222_ ), .B1(\EXU/CSRControl/_0783_ ), .B2(\EXU/CSRControl/_0149_ ), .ZN(\EXU/CSRControl/_0788_ ) );
AOI21_X1 \EXU/CSRControl/_2784_ ( .A(\EXU/CSRControl/_0788_ ), .B1(\EXU/CSRControl/_0722_ ), .B2(\EXU/CSRControl/_0750_ ), .ZN(\EXU/CSRControl/_0125_ ) );
OAI21_X1 \EXU/CSRControl/_2785_ ( .A(\EXU/CSRControl/_1222_ ), .B1(\EXU/CSRControl/_0783_ ), .B2(\EXU/CSRControl/_0150_ ), .ZN(\EXU/CSRControl/_0789_ ) );
AOI21_X1 \EXU/CSRControl/_2786_ ( .A(\EXU/CSRControl/_0789_ ), .B1(\EXU/CSRControl/_0726_ ), .B2(\EXU/CSRControl/_0750_ ), .ZN(\EXU/CSRControl/_0126_ ) );
OAI21_X1 \EXU/CSRControl/_2787_ ( .A(\EXU/CSRControl/_1222_ ), .B1(\EXU/CSRControl/_0783_ ), .B2(\EXU/CSRControl/_0151_ ), .ZN(\EXU/CSRControl/_0790_ ) );
AOI21_X1 \EXU/CSRControl/_2788_ ( .A(\EXU/CSRControl/_0790_ ), .B1(\EXU/CSRControl/_0731_ ), .B2(\EXU/CSRControl/_0750_ ), .ZN(\EXU/CSRControl/_0127_ ) );
OAI21_X1 \EXU/CSRControl/_2789_ ( .A(\EXU/CSRControl/_1222_ ), .B1(\EXU/CSRControl/_0783_ ), .B2(\EXU/CSRControl/_0152_ ), .ZN(\EXU/CSRControl/_0791_ ) );
AOI21_X1 \EXU/CSRControl/_2790_ ( .A(\EXU/CSRControl/_0791_ ), .B1(\EXU/CSRControl/_0735_ ), .B2(\EXU/CSRControl/_0750_ ), .ZN(\EXU/CSRControl/_0128_ ) );
OAI21_X1 \EXU/CSRControl/_2791_ ( .A(\EXU/CSRControl/_1222_ ), .B1(\EXU/CSRControl/_0783_ ), .B2(\EXU/CSRControl/_0153_ ), .ZN(\EXU/CSRControl/_0792_ ) );
AOI21_X1 \EXU/CSRControl/_2792_ ( .A(\EXU/CSRControl/_0792_ ), .B1(\EXU/CSRControl/_0738_ ), .B2(\EXU/CSRControl/_0750_ ), .ZN(\EXU/CSRControl/_0129_ ) );
OAI21_X1 \EXU/CSRControl/_2793_ ( .A(\EXU/CSRControl/_1222_ ), .B1(\EXU/CSRControl/_0783_ ), .B2(\EXU/CSRControl/_0155_ ), .ZN(\EXU/CSRControl/_0793_ ) );
AOI21_X1 \EXU/CSRControl/_2794_ ( .A(\EXU/CSRControl/_0793_ ), .B1(\EXU/CSRControl/_0741_ ), .B2(\EXU/CSRControl/_0750_ ), .ZN(\EXU/CSRControl/_0130_ ) );
OAI21_X1 \EXU/CSRControl/_2795_ ( .A(\EXU/CSRControl/_1222_ ), .B1(\EXU/CSRControl/_0749_ ), .B2(\EXU/CSRControl/_0156_ ), .ZN(\EXU/CSRControl/_0794_ ) );
AOI21_X1 \EXU/CSRControl/_2796_ ( .A(\EXU/CSRControl/_0794_ ), .B1(\EXU/CSRControl/_0745_ ), .B2(\EXU/CSRControl/_0750_ ), .ZN(\EXU/CSRControl/_0131_ ) );
DFF_X1 \EXU/CSRControl/_2797_ ( .D(\EXU/CSRControl/_1504_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_4_2 [3] ), .QN(\EXU/CSRControl/_1503_ ) );
DFF_X1 \EXU/CSRControl/_2798_ ( .D(\EXU/CSRControl/_1505_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_4_2 [7] ), .QN(\EXU/CSRControl/_0000_ ) );
DFF_X1 \EXU/CSRControl/_2799_ ( .D(\EXU/CSRControl/_1506_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_4_2 [11] ), .QN(\EXU/CSRControl/_1502_ ) );
DFF_X1 \EXU/CSRControl/_2800_ ( .D(\EXU/CSRControl/_1507_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_4_2 [12] ), .QN(\EXU/CSRControl/_1501_ ) );
DFF_X1 \EXU/CSRControl/_2801_ ( .D(\EXU/CSRControl/_1508_ ), .CK(clock ), .Q(\EXU/CSRControl/priv [0] ), .QN(\EXU/CSRControl/_1500_ ) );
DFF_X1 \EXU/CSRControl/_2802_ ( .D(\EXU/CSRControl/_1509_ ), .CK(clock ), .Q(\EXU/CSRControl/priv [1] ), .QN(\EXU/CSRControl/_1499_ ) );
DFF_X1 \EXU/CSRControl/_2803_ ( .D(\EXU/CSRControl/_1510_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_4_2 [0] ), .QN(\EXU/CSRControl/_1498_ ) );
DFF_X1 \EXU/CSRControl/_2804_ ( .D(\EXU/CSRControl/_1511_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_4_2 [1] ), .QN(\EXU/CSRControl/_1497_ ) );
DFF_X1 \EXU/CSRControl/_2805_ ( .D(\EXU/CSRControl/_1512_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_4_2 [2] ), .QN(\EXU/CSRControl/_1496_ ) );
DFF_X1 \EXU/CSRControl/_2806_ ( .D(\EXU/CSRControl/_1513_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_4_2 [4] ), .QN(\EXU/CSRControl/_1495_ ) );
DFF_X1 \EXU/CSRControl/_2807_ ( .D(\EXU/CSRControl/_1514_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_4_2 [5] ), .QN(\EXU/CSRControl/_1494_ ) );
DFF_X1 \EXU/CSRControl/_2808_ ( .D(\EXU/CSRControl/_1515_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_4_2 [6] ), .QN(\EXU/CSRControl/_1493_ ) );
DFF_X1 \EXU/CSRControl/_2809_ ( .D(\EXU/CSRControl/_1516_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_4_2 [8] ), .QN(\EXU/CSRControl/_1492_ ) );
DFF_X1 \EXU/CSRControl/_2810_ ( .D(\EXU/CSRControl/_1517_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_4_2 [9] ), .QN(\EXU/CSRControl/_1491_ ) );
DFF_X1 \EXU/CSRControl/_2811_ ( .D(\EXU/CSRControl/_1518_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_4_2 [10] ), .QN(\EXU/CSRControl/_1490_ ) );
DFF_X1 \EXU/CSRControl/_2812_ ( .D(\EXU/CSRControl/_1519_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_4_2 [13] ), .QN(\EXU/CSRControl/_1489_ ) );
DFF_X1 \EXU/CSRControl/_2813_ ( .D(\EXU/CSRControl/_1520_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_4_2 [14] ), .QN(\EXU/CSRControl/_1488_ ) );
DFF_X1 \EXU/CSRControl/_2814_ ( .D(\EXU/CSRControl/_1521_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_4_2 [15] ), .QN(\EXU/CSRControl/_1487_ ) );
DFF_X1 \EXU/CSRControl/_2815_ ( .D(\EXU/CSRControl/_1522_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_4_2 [16] ), .QN(\EXU/CSRControl/_1486_ ) );
DFF_X1 \EXU/CSRControl/_2816_ ( .D(\EXU/CSRControl/_1523_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_4_2 [17] ), .QN(\EXU/CSRControl/_1485_ ) );
DFF_X1 \EXU/CSRControl/_2817_ ( .D(\EXU/CSRControl/_1524_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_4_2 [18] ), .QN(\EXU/CSRControl/_1484_ ) );
DFF_X1 \EXU/CSRControl/_2818_ ( .D(\EXU/CSRControl/_1525_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_4_2 [19] ), .QN(\EXU/CSRControl/_1483_ ) );
DFF_X1 \EXU/CSRControl/_2819_ ( .D(\EXU/CSRControl/_1526_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_4_2 [20] ), .QN(\EXU/CSRControl/_1482_ ) );
DFF_X1 \EXU/CSRControl/_2820_ ( .D(\EXU/CSRControl/_1527_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_4_2 [21] ), .QN(\EXU/CSRControl/_1481_ ) );
DFF_X1 \EXU/CSRControl/_2821_ ( .D(\EXU/CSRControl/_1528_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_4_2 [22] ), .QN(\EXU/CSRControl/_1480_ ) );
DFF_X1 \EXU/CSRControl/_2822_ ( .D(\EXU/CSRControl/_1529_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_4_2 [23] ), .QN(\EXU/CSRControl/_1479_ ) );
DFF_X1 \EXU/CSRControl/_2823_ ( .D(\EXU/CSRControl/_1530_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_4_2 [24] ), .QN(\EXU/CSRControl/_1478_ ) );
DFF_X1 \EXU/CSRControl/_2824_ ( .D(\EXU/CSRControl/_1531_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_4_2 [25] ), .QN(\EXU/CSRControl/_1477_ ) );
DFF_X1 \EXU/CSRControl/_2825_ ( .D(\EXU/CSRControl/_1532_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_4_2 [26] ), .QN(\EXU/CSRControl/_1476_ ) );
DFF_X1 \EXU/CSRControl/_2826_ ( .D(\EXU/CSRControl/_1533_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_4_2 [27] ), .QN(\EXU/CSRControl/_1475_ ) );
DFF_X1 \EXU/CSRControl/_2827_ ( .D(\EXU/CSRControl/_1534_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_4_2 [28] ), .QN(\EXU/CSRControl/_1474_ ) );
DFF_X1 \EXU/CSRControl/_2828_ ( .D(\EXU/CSRControl/_1535_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_4_2 [29] ), .QN(\EXU/CSRControl/_1473_ ) );
DFF_X1 \EXU/CSRControl/_2829_ ( .D(\EXU/CSRControl/_1536_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_4_2 [30] ), .QN(\EXU/CSRControl/_1472_ ) );
DFF_X1 \EXU/CSRControl/_2830_ ( .D(\EXU/CSRControl/_1537_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_4_2 [31] ), .QN(\EXU/CSRControl/_1471_ ) );
DFF_X1 \EXU/CSRControl/_2831_ ( .D(\EXU/CSRControl/_1538_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_2_2 [0] ), .QN(\EXU/CSRControl/_1470_ ) );
DFF_X1 \EXU/CSRControl/_2832_ ( .D(\EXU/CSRControl/_1539_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_2_2 [1] ), .QN(\EXU/CSRControl/_1469_ ) );
DFF_X1 \EXU/CSRControl/_2833_ ( .D(\EXU/CSRControl/_1540_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_2_2 [2] ), .QN(\EXU/CSRControl/_1468_ ) );
DFF_X1 \EXU/CSRControl/_2834_ ( .D(\EXU/CSRControl/_1541_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_2_2 [3] ), .QN(\EXU/CSRControl/_1467_ ) );
DFF_X1 \EXU/CSRControl/_2835_ ( .D(\EXU/CSRControl/_1542_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_2_2 [4] ), .QN(\EXU/CSRControl/_1466_ ) );
DFF_X1 \EXU/CSRControl/_2836_ ( .D(\EXU/CSRControl/_1543_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_2_2 [5] ), .QN(\EXU/CSRControl/_1465_ ) );
DFF_X1 \EXU/CSRControl/_2837_ ( .D(\EXU/CSRControl/_1544_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_2_2 [6] ), .QN(\EXU/CSRControl/_1464_ ) );
DFF_X1 \EXU/CSRControl/_2838_ ( .D(\EXU/CSRControl/_1545_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_2_2 [7] ), .QN(\EXU/CSRControl/_1463_ ) );
DFF_X1 \EXU/CSRControl/_2839_ ( .D(\EXU/CSRControl/_1546_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_2_2 [8] ), .QN(\EXU/CSRControl/_1462_ ) );
DFF_X1 \EXU/CSRControl/_2840_ ( .D(\EXU/CSRControl/_1547_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_2_2 [9] ), .QN(\EXU/CSRControl/_1461_ ) );
DFF_X1 \EXU/CSRControl/_2841_ ( .D(\EXU/CSRControl/_1548_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_2_2 [10] ), .QN(\EXU/CSRControl/_1460_ ) );
DFF_X1 \EXU/CSRControl/_2842_ ( .D(\EXU/CSRControl/_1549_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_2_2 [11] ), .QN(\EXU/CSRControl/_1459_ ) );
DFF_X1 \EXU/CSRControl/_2843_ ( .D(\EXU/CSRControl/_1550_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_2_2 [12] ), .QN(\EXU/CSRControl/_1458_ ) );
DFF_X1 \EXU/CSRControl/_2844_ ( .D(\EXU/CSRControl/_1551_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_2_2 [13] ), .QN(\EXU/CSRControl/_1457_ ) );
DFF_X1 \EXU/CSRControl/_2845_ ( .D(\EXU/CSRControl/_1552_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_2_2 [14] ), .QN(\EXU/CSRControl/_1456_ ) );
DFF_X1 \EXU/CSRControl/_2846_ ( .D(\EXU/CSRControl/_1553_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_2_2 [15] ), .QN(\EXU/CSRControl/_1455_ ) );
DFF_X1 \EXU/CSRControl/_2847_ ( .D(\EXU/CSRControl/_1554_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_2_2 [16] ), .QN(\EXU/CSRControl/_1454_ ) );
DFF_X1 \EXU/CSRControl/_2848_ ( .D(\EXU/CSRControl/_1555_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_2_2 [17] ), .QN(\EXU/CSRControl/_1453_ ) );
DFF_X1 \EXU/CSRControl/_2849_ ( .D(\EXU/CSRControl/_1556_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_2_2 [18] ), .QN(\EXU/CSRControl/_1452_ ) );
DFF_X1 \EXU/CSRControl/_2850_ ( .D(\EXU/CSRControl/_1557_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_2_2 [19] ), .QN(\EXU/CSRControl/_1451_ ) );
DFF_X1 \EXU/CSRControl/_2851_ ( .D(\EXU/CSRControl/_1558_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_2_2 [20] ), .QN(\EXU/CSRControl/_1450_ ) );
DFF_X1 \EXU/CSRControl/_2852_ ( .D(\EXU/CSRControl/_1559_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_2_2 [21] ), .QN(\EXU/CSRControl/_1449_ ) );
DFF_X1 \EXU/CSRControl/_2853_ ( .D(\EXU/CSRControl/_1560_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_2_2 [22] ), .QN(\EXU/CSRControl/_1448_ ) );
DFF_X1 \EXU/CSRControl/_2854_ ( .D(\EXU/CSRControl/_1561_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_2_2 [23] ), .QN(\EXU/CSRControl/_1447_ ) );
DFF_X1 \EXU/CSRControl/_2855_ ( .D(\EXU/CSRControl/_1562_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_2_2 [24] ), .QN(\EXU/CSRControl/_1446_ ) );
DFF_X1 \EXU/CSRControl/_2856_ ( .D(\EXU/CSRControl/_1563_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_2_2 [25] ), .QN(\EXU/CSRControl/_1445_ ) );
DFF_X1 \EXU/CSRControl/_2857_ ( .D(\EXU/CSRControl/_1564_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_2_2 [26] ), .QN(\EXU/CSRControl/_1444_ ) );
DFF_X1 \EXU/CSRControl/_2858_ ( .D(\EXU/CSRControl/_1565_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_2_2 [27] ), .QN(\EXU/CSRControl/_1443_ ) );
DFF_X1 \EXU/CSRControl/_2859_ ( .D(\EXU/CSRControl/_1566_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_2_2 [28] ), .QN(\EXU/CSRControl/_1442_ ) );
DFF_X1 \EXU/CSRControl/_2860_ ( .D(\EXU/CSRControl/_1567_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_2_2 [29] ), .QN(\EXU/CSRControl/_1441_ ) );
DFF_X1 \EXU/CSRControl/_2861_ ( .D(\EXU/CSRControl/_1568_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_2_2 [30] ), .QN(\EXU/CSRControl/_1440_ ) );
DFF_X1 \EXU/CSRControl/_2862_ ( .D(\EXU/CSRControl/_1569_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_2_2 [31] ), .QN(\EXU/CSRControl/_1439_ ) );
DFF_X1 \EXU/CSRControl/_2863_ ( .D(\EXU/CSRControl/_1570_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_3_2 [0] ), .QN(\EXU/CSRControl/_1438_ ) );
DFF_X1 \EXU/CSRControl/_2864_ ( .D(\EXU/CSRControl/_1571_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_3_2 [1] ), .QN(\EXU/CSRControl/_1437_ ) );
DFF_X1 \EXU/CSRControl/_2865_ ( .D(\EXU/CSRControl/_1572_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_3_2 [2] ), .QN(\EXU/CSRControl/_1436_ ) );
DFF_X1 \EXU/CSRControl/_2866_ ( .D(\EXU/CSRControl/_1573_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_3_2 [3] ), .QN(\EXU/CSRControl/_1435_ ) );
DFF_X1 \EXU/CSRControl/_2867_ ( .D(\EXU/CSRControl/_1574_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_3_2 [4] ), .QN(\EXU/CSRControl/_1434_ ) );
DFF_X1 \EXU/CSRControl/_2868_ ( .D(\EXU/CSRControl/_1575_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_3_2 [5] ), .QN(\EXU/CSRControl/_1433_ ) );
DFF_X1 \EXU/CSRControl/_2869_ ( .D(\EXU/CSRControl/_1576_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_3_2 [6] ), .QN(\EXU/CSRControl/_1432_ ) );
DFF_X1 \EXU/CSRControl/_2870_ ( .D(\EXU/CSRControl/_1577_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_3_2 [7] ), .QN(\EXU/CSRControl/_1431_ ) );
DFF_X1 \EXU/CSRControl/_2871_ ( .D(\EXU/CSRControl/_1578_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_3_2 [8] ), .QN(\EXU/CSRControl/_1430_ ) );
DFF_X1 \EXU/CSRControl/_2872_ ( .D(\EXU/CSRControl/_1579_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_3_2 [9] ), .QN(\EXU/CSRControl/_1429_ ) );
DFF_X1 \EXU/CSRControl/_2873_ ( .D(\EXU/CSRControl/_1580_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_3_2 [10] ), .QN(\EXU/CSRControl/_1428_ ) );
DFF_X1 \EXU/CSRControl/_2874_ ( .D(\EXU/CSRControl/_1581_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_3_2 [11] ), .QN(\EXU/CSRControl/_1427_ ) );
DFF_X1 \EXU/CSRControl/_2875_ ( .D(\EXU/CSRControl/_1582_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_3_2 [12] ), .QN(\EXU/CSRControl/_1426_ ) );
DFF_X1 \EXU/CSRControl/_2876_ ( .D(\EXU/CSRControl/_1583_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_3_2 [13] ), .QN(\EXU/CSRControl/_1425_ ) );
DFF_X1 \EXU/CSRControl/_2877_ ( .D(\EXU/CSRControl/_1584_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_3_2 [14] ), .QN(\EXU/CSRControl/_1424_ ) );
DFF_X1 \EXU/CSRControl/_2878_ ( .D(\EXU/CSRControl/_1585_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_3_2 [15] ), .QN(\EXU/CSRControl/_1423_ ) );
DFF_X1 \EXU/CSRControl/_2879_ ( .D(\EXU/CSRControl/_1586_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_3_2 [16] ), .QN(\EXU/CSRControl/_1422_ ) );
DFF_X1 \EXU/CSRControl/_2880_ ( .D(\EXU/CSRControl/_1587_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_3_2 [17] ), .QN(\EXU/CSRControl/_1421_ ) );
DFF_X1 \EXU/CSRControl/_2881_ ( .D(\EXU/CSRControl/_1588_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_3_2 [18] ), .QN(\EXU/CSRControl/_1420_ ) );
DFF_X1 \EXU/CSRControl/_2882_ ( .D(\EXU/CSRControl/_1589_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_3_2 [19] ), .QN(\EXU/CSRControl/_1419_ ) );
DFF_X1 \EXU/CSRControl/_2883_ ( .D(\EXU/CSRControl/_1590_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_3_2 [20] ), .QN(\EXU/CSRControl/_1418_ ) );
DFF_X1 \EXU/CSRControl/_2884_ ( .D(\EXU/CSRControl/_1591_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_3_2 [21] ), .QN(\EXU/CSRControl/_1417_ ) );
DFF_X1 \EXU/CSRControl/_2885_ ( .D(\EXU/CSRControl/_1592_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_3_2 [22] ), .QN(\EXU/CSRControl/_1416_ ) );
DFF_X1 \EXU/CSRControl/_2886_ ( .D(\EXU/CSRControl/_1593_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_3_2 [23] ), .QN(\EXU/CSRControl/_1415_ ) );
DFF_X1 \EXU/CSRControl/_2887_ ( .D(\EXU/CSRControl/_1594_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_3_2 [24] ), .QN(\EXU/CSRControl/_1414_ ) );
DFF_X1 \EXU/CSRControl/_2888_ ( .D(\EXU/CSRControl/_1595_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_3_2 [25] ), .QN(\EXU/CSRControl/_1413_ ) );
DFF_X1 \EXU/CSRControl/_2889_ ( .D(\EXU/CSRControl/_1596_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_3_2 [26] ), .QN(\EXU/CSRControl/_1412_ ) );
DFF_X1 \EXU/CSRControl/_2890_ ( .D(\EXU/CSRControl/_1597_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_3_2 [27] ), .QN(\EXU/CSRControl/_1411_ ) );
DFF_X1 \EXU/CSRControl/_2891_ ( .D(\EXU/CSRControl/_1598_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_3_2 [28] ), .QN(\EXU/CSRControl/_1410_ ) );
DFF_X1 \EXU/CSRControl/_2892_ ( .D(\EXU/CSRControl/_1599_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_3_2 [29] ), .QN(\EXU/CSRControl/_1409_ ) );
DFF_X1 \EXU/CSRControl/_2893_ ( .D(\EXU/CSRControl/_1600_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_3_2 [30] ), .QN(\EXU/CSRControl/_1408_ ) );
DFF_X1 \EXU/CSRControl/_2894_ ( .D(\EXU/CSRControl/_1601_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_3_2 [31] ), .QN(\EXU/CSRControl/_1407_ ) );
DFF_X1 \EXU/CSRControl/_2895_ ( .D(\EXU/CSRControl/_1602_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_0_2 [0] ), .QN(\EXU/CSRControl/_1406_ ) );
DFF_X1 \EXU/CSRControl/_2896_ ( .D(\EXU/CSRControl/_1603_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_0_2 [1] ), .QN(\EXU/CSRControl/_1405_ ) );
DFF_X1 \EXU/CSRControl/_2897_ ( .D(\EXU/CSRControl/_1604_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_0_2 [2] ), .QN(\EXU/CSRControl/_1404_ ) );
DFF_X1 \EXU/CSRControl/_2898_ ( .D(\EXU/CSRControl/_1605_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_0_2 [3] ), .QN(\EXU/CSRControl/_1403_ ) );
DFF_X1 \EXU/CSRControl/_2899_ ( .D(\EXU/CSRControl/_1606_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_0_2 [4] ), .QN(\EXU/CSRControl/_1402_ ) );
DFF_X1 \EXU/CSRControl/_2900_ ( .D(\EXU/CSRControl/_1607_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_0_2 [5] ), .QN(\EXU/CSRControl/_1401_ ) );
DFF_X1 \EXU/CSRControl/_2901_ ( .D(\EXU/CSRControl/_1608_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_0_2 [6] ), .QN(\EXU/CSRControl/_1400_ ) );
DFF_X1 \EXU/CSRControl/_2902_ ( .D(\EXU/CSRControl/_1609_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_0_2 [7] ), .QN(\EXU/CSRControl/_1399_ ) );
DFF_X1 \EXU/CSRControl/_2903_ ( .D(\EXU/CSRControl/_1610_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_0_2 [8] ), .QN(\EXU/CSRControl/_1398_ ) );
DFF_X1 \EXU/CSRControl/_2904_ ( .D(\EXU/CSRControl/_1611_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_0_2 [9] ), .QN(\EXU/CSRControl/_1397_ ) );
DFF_X1 \EXU/CSRControl/_2905_ ( .D(\EXU/CSRControl/_1612_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_0_2 [10] ), .QN(\EXU/CSRControl/_1396_ ) );
DFF_X1 \EXU/CSRControl/_2906_ ( .D(\EXU/CSRControl/_1613_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_0_2 [11] ), .QN(\EXU/CSRControl/_1395_ ) );
DFF_X1 \EXU/CSRControl/_2907_ ( .D(\EXU/CSRControl/_1614_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_0_2 [12] ), .QN(\EXU/CSRControl/_1394_ ) );
DFF_X1 \EXU/CSRControl/_2908_ ( .D(\EXU/CSRControl/_1615_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_0_2 [13] ), .QN(\EXU/CSRControl/_1393_ ) );
DFF_X1 \EXU/CSRControl/_2909_ ( .D(\EXU/CSRControl/_1616_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_0_2 [14] ), .QN(\EXU/CSRControl/_1392_ ) );
DFF_X1 \EXU/CSRControl/_2910_ ( .D(\EXU/CSRControl/_1617_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_0_2 [15] ), .QN(\EXU/CSRControl/_1391_ ) );
DFF_X1 \EXU/CSRControl/_2911_ ( .D(\EXU/CSRControl/_1618_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_0_2 [16] ), .QN(\EXU/CSRControl/_1390_ ) );
DFF_X1 \EXU/CSRControl/_2912_ ( .D(\EXU/CSRControl/_1619_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_0_2 [17] ), .QN(\EXU/CSRControl/_1389_ ) );
DFF_X1 \EXU/CSRControl/_2913_ ( .D(\EXU/CSRControl/_1620_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_0_2 [18] ), .QN(\EXU/CSRControl/_1388_ ) );
DFF_X1 \EXU/CSRControl/_2914_ ( .D(\EXU/CSRControl/_1621_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_0_2 [19] ), .QN(\EXU/CSRControl/_1387_ ) );
DFF_X1 \EXU/CSRControl/_2915_ ( .D(\EXU/CSRControl/_1622_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_0_2 [20] ), .QN(\EXU/CSRControl/_1386_ ) );
DFF_X1 \EXU/CSRControl/_2916_ ( .D(\EXU/CSRControl/_1623_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_0_2 [21] ), .QN(\EXU/CSRControl/_1385_ ) );
DFF_X1 \EXU/CSRControl/_2917_ ( .D(\EXU/CSRControl/_1624_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_0_2 [22] ), .QN(\EXU/CSRControl/_1384_ ) );
DFF_X1 \EXU/CSRControl/_2918_ ( .D(\EXU/CSRControl/_1625_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_0_2 [23] ), .QN(\EXU/CSRControl/_1383_ ) );
DFF_X1 \EXU/CSRControl/_2919_ ( .D(\EXU/CSRControl/_1626_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_0_2 [24] ), .QN(\EXU/CSRControl/_1382_ ) );
DFF_X1 \EXU/CSRControl/_2920_ ( .D(\EXU/CSRControl/_1627_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_0_2 [25] ), .QN(\EXU/CSRControl/_1381_ ) );
DFF_X1 \EXU/CSRControl/_2921_ ( .D(\EXU/CSRControl/_1628_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_0_2 [26] ), .QN(\EXU/CSRControl/_1380_ ) );
DFF_X1 \EXU/CSRControl/_2922_ ( .D(\EXU/CSRControl/_1629_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_0_2 [27] ), .QN(\EXU/CSRControl/_1379_ ) );
DFF_X1 \EXU/CSRControl/_2923_ ( .D(\EXU/CSRControl/_1630_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_0_2 [28] ), .QN(\EXU/CSRControl/_1378_ ) );
DFF_X1 \EXU/CSRControl/_2924_ ( .D(\EXU/CSRControl/_1631_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_0_2 [29] ), .QN(\EXU/CSRControl/_1377_ ) );
DFF_X1 \EXU/CSRControl/_2925_ ( .D(\EXU/CSRControl/_1632_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_0_2 [30] ), .QN(\EXU/CSRControl/_1376_ ) );
DFF_X1 \EXU/CSRControl/_2926_ ( .D(\EXU/CSRControl/_1633_ ), .CK(clock ), .Q(\EXU/CSRControl/csrs_0_2 [31] ), .QN(\EXU/CSRControl/_1375_ ) );
BUF_X1 \EXU/CSRControl/_2927_ ( .A(\EXU/in_imm [1] ), .Z(\EXU/CSRControl/_0263_ ) );
BUF_X1 \EXU/CSRControl/_2928_ ( .A(\EXU/in_imm [0] ), .Z(\EXU/CSRControl/_0260_ ) );
BUF_X1 \EXU/CSRControl/_2929_ ( .A(\EXU/in_imm [3] ), .Z(\EXU/CSRControl/_0265_ ) );
BUF_X1 \EXU/CSRControl/_2930_ ( .A(\EXU/in_imm [2] ), .Z(\EXU/CSRControl/_0264_ ) );
BUF_X1 \EXU/CSRControl/_2931_ ( .A(\EXU/in_imm [5] ), .Z(\EXU/CSRControl/_0267_ ) );
BUF_X1 \EXU/CSRControl/_2932_ ( .A(\EXU/in_imm [4] ), .Z(\EXU/CSRControl/_0266_ ) );
BUF_X1 \EXU/CSRControl/_2933_ ( .A(\EXU/in_imm [7] ), .Z(\EXU/CSRControl/_0269_ ) );
BUF_X1 \EXU/CSRControl/_2934_ ( .A(\EXU/in_imm [6] ), .Z(\EXU/CSRControl/_0268_ ) );
BUF_X1 \EXU/CSRControl/_2935_ ( .A(\EXU/in_imm [9] ), .Z(\EXU/CSRControl/_0271_ ) );
BUF_X1 \EXU/CSRControl/_2936_ ( .A(\EXU/in_imm [8] ), .Z(\EXU/CSRControl/_0270_ ) );
BUF_X1 \EXU/CSRControl/_2937_ ( .A(\EXU/_0033_ ), .Z(\EXU/CSRControl/_0273_ ) );
BUF_X1 \EXU/CSRControl/_2938_ ( .A(\EXU/_0032_ ), .Z(\EXU/CSRControl/_0272_ ) );
BUF_X1 \EXU/CSRControl/_2939_ ( .A(\EXU/_0034_ ), .Z(\EXU/CSRControl/_0274_ ) );
BUF_X1 \EXU/CSRControl/_2940_ ( .A(reset ), .Z(\EXU/CSRControl/_1374_ ) );
BUF_X1 \EXU/CSRControl/_2941_ ( .A(\EXU/CSRControl/csrs_4_2 [0] ), .Z(\EXU/CSRControl/_0228_ ) );
BUF_X1 \EXU/CSRControl/_2942_ ( .A(\EXU/CSRControl/csrs_3_2 [0] ), .Z(\EXU/CSRControl/_0196_ ) );
BUF_X1 \EXU/CSRControl/_2943_ ( .A(\EXU/CSRControl/csrs_2_2 [0] ), .Z(\EXU/CSRControl/_0164_ ) );
BUF_X1 \EXU/CSRControl/_2944_ ( .A(\EXU/in_imm [11] ), .Z(\EXU/CSRControl/_0262_ ) );
BUF_X1 \EXU/CSRControl/_2945_ ( .A(\EXU/in_imm [10] ), .Z(\EXU/CSRControl/_0261_ ) );
BUF_X1 \EXU/CSRControl/_2946_ ( .A(\EXU/CSRControl/csrs_0_2 [0] ), .Z(\EXU/CSRControl/_0132_ ) );
BUF_X1 \EXU/CSRControl/_2947_ ( .A(\EXU/CSRControl/_0307_ ), .Z(\_EXU_io_out_bits_csrOut [0] ) );
BUF_X1 \EXU/CSRControl/_2948_ ( .A(\EXU/CSRControl/csrs_4_2 [1] ), .Z(\EXU/CSRControl/_0239_ ) );
BUF_X1 \EXU/CSRControl/_2949_ ( .A(\EXU/CSRControl/csrs_3_2 [1] ), .Z(\EXU/CSRControl/_0207_ ) );
BUF_X1 \EXU/CSRControl/_2950_ ( .A(\EXU/CSRControl/csrs_2_2 [1] ), .Z(\EXU/CSRControl/_0175_ ) );
BUF_X1 \EXU/CSRControl/_2951_ ( .A(\EXU/CSRControl/csrs_0_2 [1] ), .Z(\EXU/CSRControl/_0143_ ) );
BUF_X1 \EXU/CSRControl/_2952_ ( .A(\EXU/CSRControl/_0318_ ), .Z(\_EXU_io_out_bits_csrOut [1] ) );
BUF_X1 \EXU/CSRControl/_2953_ ( .A(\EXU/CSRControl/csrs_4_2 [2] ), .Z(\EXU/CSRControl/_0250_ ) );
BUF_X1 \EXU/CSRControl/_2954_ ( .A(\EXU/CSRControl/csrs_3_2 [2] ), .Z(\EXU/CSRControl/_0218_ ) );
BUF_X1 \EXU/CSRControl/_2955_ ( .A(\EXU/CSRControl/csrs_2_2 [2] ), .Z(\EXU/CSRControl/_0186_ ) );
BUF_X1 \EXU/CSRControl/_2956_ ( .A(\EXU/CSRControl/csrs_0_2 [2] ), .Z(\EXU/CSRControl/_0154_ ) );
BUF_X1 \EXU/CSRControl/_2957_ ( .A(\EXU/CSRControl/_0329_ ), .Z(\_EXU_io_out_bits_csrOut [2] ) );
BUF_X1 \EXU/CSRControl/_2958_ ( .A(\EXU/CSRControl/csrs_4_2 [3] ), .Z(\EXU/CSRControl/_0253_ ) );
BUF_X1 \EXU/CSRControl/_2959_ ( .A(\EXU/CSRControl/csrs_3_2 [3] ), .Z(\EXU/CSRControl/_0221_ ) );
BUF_X1 \EXU/CSRControl/_2960_ ( .A(\EXU/CSRControl/csrs_2_2 [3] ), .Z(\EXU/CSRControl/_0189_ ) );
BUF_X1 \EXU/CSRControl/_2961_ ( .A(\EXU/CSRControl/csrs_0_2 [3] ), .Z(\EXU/CSRControl/_0157_ ) );
BUF_X1 \EXU/CSRControl/_2962_ ( .A(\EXU/CSRControl/_0332_ ), .Z(\_EXU_io_out_bits_csrOut [3] ) );
BUF_X1 \EXU/CSRControl/_2963_ ( .A(\EXU/CSRControl/csrs_4_2 [4] ), .Z(\EXU/CSRControl/_0254_ ) );
BUF_X1 \EXU/CSRControl/_2964_ ( .A(\EXU/CSRControl/csrs_3_2 [4] ), .Z(\EXU/CSRControl/_0222_ ) );
BUF_X1 \EXU/CSRControl/_2965_ ( .A(\EXU/CSRControl/csrs_2_2 [4] ), .Z(\EXU/CSRControl/_0190_ ) );
BUF_X1 \EXU/CSRControl/_2966_ ( .A(\EXU/CSRControl/csrs_0_2 [4] ), .Z(\EXU/CSRControl/_0158_ ) );
BUF_X1 \EXU/CSRControl/_2967_ ( .A(\EXU/CSRControl/_0333_ ), .Z(\_EXU_io_out_bits_csrOut [4] ) );
BUF_X1 \EXU/CSRControl/_2968_ ( .A(\EXU/CSRControl/csrs_4_2 [5] ), .Z(\EXU/CSRControl/_0255_ ) );
BUF_X1 \EXU/CSRControl/_2969_ ( .A(\EXU/CSRControl/csrs_3_2 [5] ), .Z(\EXU/CSRControl/_0223_ ) );
BUF_X1 \EXU/CSRControl/_2970_ ( .A(\EXU/CSRControl/csrs_2_2 [5] ), .Z(\EXU/CSRControl/_0191_ ) );
BUF_X1 \EXU/CSRControl/_2971_ ( .A(\EXU/CSRControl/csrs_0_2 [5] ), .Z(\EXU/CSRControl/_0159_ ) );
BUF_X1 \EXU/CSRControl/_2972_ ( .A(\EXU/CSRControl/_0334_ ), .Z(\_EXU_io_out_bits_csrOut [5] ) );
BUF_X1 \EXU/CSRControl/_2973_ ( .A(\EXU/CSRControl/csrs_4_2 [6] ), .Z(\EXU/CSRControl/_0256_ ) );
BUF_X1 \EXU/CSRControl/_2974_ ( .A(\EXU/CSRControl/csrs_3_2 [6] ), .Z(\EXU/CSRControl/_0224_ ) );
BUF_X1 \EXU/CSRControl/_2975_ ( .A(\EXU/CSRControl/csrs_2_2 [6] ), .Z(\EXU/CSRControl/_0192_ ) );
BUF_X1 \EXU/CSRControl/_2976_ ( .A(\EXU/CSRControl/csrs_0_2 [6] ), .Z(\EXU/CSRControl/_0160_ ) );
BUF_X1 \EXU/CSRControl/_2977_ ( .A(\EXU/CSRControl/_0335_ ), .Z(\_EXU_io_out_bits_csrOut [6] ) );
BUF_X1 \EXU/CSRControl/_2978_ ( .A(\EXU/CSRControl/csrs_4_2 [7] ), .Z(\EXU/CSRControl/_0257_ ) );
BUF_X1 \EXU/CSRControl/_2979_ ( .A(\EXU/CSRControl/csrs_3_2 [7] ), .Z(\EXU/CSRControl/_0225_ ) );
BUF_X1 \EXU/CSRControl/_2980_ ( .A(\EXU/CSRControl/csrs_2_2 [7] ), .Z(\EXU/CSRControl/_0193_ ) );
BUF_X1 \EXU/CSRControl/_2981_ ( .A(\EXU/CSRControl/csrs_0_2 [7] ), .Z(\EXU/CSRControl/_0161_ ) );
BUF_X1 \EXU/CSRControl/_2982_ ( .A(\EXU/CSRControl/_0336_ ), .Z(\_EXU_io_out_bits_csrOut [7] ) );
BUF_X1 \EXU/CSRControl/_2983_ ( .A(\EXU/CSRControl/csrs_4_2 [8] ), .Z(\EXU/CSRControl/_0258_ ) );
BUF_X1 \EXU/CSRControl/_2984_ ( .A(\EXU/CSRControl/csrs_3_2 [8] ), .Z(\EXU/CSRControl/_0226_ ) );
BUF_X1 \EXU/CSRControl/_2985_ ( .A(\EXU/CSRControl/csrs_2_2 [8] ), .Z(\EXU/CSRControl/_0194_ ) );
BUF_X1 \EXU/CSRControl/_2986_ ( .A(\EXU/CSRControl/csrs_0_2 [8] ), .Z(\EXU/CSRControl/_0162_ ) );
BUF_X1 \EXU/CSRControl/_2987_ ( .A(\EXU/CSRControl/_0337_ ), .Z(\_EXU_io_out_bits_csrOut [8] ) );
BUF_X1 \EXU/CSRControl/_2988_ ( .A(\EXU/CSRControl/csrs_4_2 [9] ), .Z(\EXU/CSRControl/_0259_ ) );
BUF_X1 \EXU/CSRControl/_2989_ ( .A(\EXU/CSRControl/csrs_3_2 [9] ), .Z(\EXU/CSRControl/_0227_ ) );
BUF_X1 \EXU/CSRControl/_2990_ ( .A(\EXU/CSRControl/csrs_2_2 [9] ), .Z(\EXU/CSRControl/_0195_ ) );
BUF_X1 \EXU/CSRControl/_2991_ ( .A(\EXU/CSRControl/csrs_0_2 [9] ), .Z(\EXU/CSRControl/_0163_ ) );
BUF_X1 \EXU/CSRControl/_2992_ ( .A(\EXU/CSRControl/_0338_ ), .Z(\_EXU_io_out_bits_csrOut [9] ) );
BUF_X1 \EXU/CSRControl/_2993_ ( .A(\EXU/CSRControl/csrs_4_2 [10] ), .Z(\EXU/CSRControl/_0229_ ) );
BUF_X1 \EXU/CSRControl/_2994_ ( .A(\EXU/CSRControl/csrs_3_2 [10] ), .Z(\EXU/CSRControl/_0197_ ) );
BUF_X1 \EXU/CSRControl/_2995_ ( .A(\EXU/CSRControl/csrs_2_2 [10] ), .Z(\EXU/CSRControl/_0165_ ) );
BUF_X1 \EXU/CSRControl/_2996_ ( .A(\EXU/CSRControl/csrs_0_2 [10] ), .Z(\EXU/CSRControl/_0133_ ) );
BUF_X1 \EXU/CSRControl/_2997_ ( .A(\EXU/CSRControl/_0308_ ), .Z(\_EXU_io_out_bits_csrOut [10] ) );
BUF_X1 \EXU/CSRControl/_2998_ ( .A(\EXU/CSRControl/csrs_4_2 [11] ), .Z(\EXU/CSRControl/_0230_ ) );
BUF_X1 \EXU/CSRControl/_2999_ ( .A(\EXU/CSRControl/csrs_3_2 [11] ), .Z(\EXU/CSRControl/_0198_ ) );
BUF_X1 \EXU/CSRControl/_3000_ ( .A(\EXU/CSRControl/csrs_2_2 [11] ), .Z(\EXU/CSRControl/_0166_ ) );
BUF_X1 \EXU/CSRControl/_3001_ ( .A(\EXU/CSRControl/csrs_0_2 [11] ), .Z(\EXU/CSRControl/_0134_ ) );
BUF_X1 \EXU/CSRControl/_3002_ ( .A(\EXU/CSRControl/_0309_ ), .Z(\_EXU_io_out_bits_csrOut [11] ) );
BUF_X1 \EXU/CSRControl/_3003_ ( .A(\EXU/CSRControl/csrs_4_2 [12] ), .Z(\EXU/CSRControl/_0231_ ) );
BUF_X1 \EXU/CSRControl/_3004_ ( .A(\EXU/CSRControl/csrs_3_2 [12] ), .Z(\EXU/CSRControl/_0199_ ) );
BUF_X1 \EXU/CSRControl/_3005_ ( .A(\EXU/CSRControl/csrs_2_2 [12] ), .Z(\EXU/CSRControl/_0167_ ) );
BUF_X1 \EXU/CSRControl/_3006_ ( .A(\EXU/CSRControl/csrs_0_2 [12] ), .Z(\EXU/CSRControl/_0135_ ) );
BUF_X1 \EXU/CSRControl/_3007_ ( .A(\EXU/CSRControl/_0310_ ), .Z(\_EXU_io_out_bits_csrOut [12] ) );
BUF_X1 \EXU/CSRControl/_3008_ ( .A(\EXU/CSRControl/csrs_4_2 [13] ), .Z(\EXU/CSRControl/_0232_ ) );
BUF_X1 \EXU/CSRControl/_3009_ ( .A(\EXU/CSRControl/csrs_3_2 [13] ), .Z(\EXU/CSRControl/_0200_ ) );
BUF_X1 \EXU/CSRControl/_3010_ ( .A(\EXU/CSRControl/csrs_2_2 [13] ), .Z(\EXU/CSRControl/_0168_ ) );
BUF_X1 \EXU/CSRControl/_3011_ ( .A(\EXU/CSRControl/csrs_0_2 [13] ), .Z(\EXU/CSRControl/_0136_ ) );
BUF_X1 \EXU/CSRControl/_3012_ ( .A(\EXU/CSRControl/_0311_ ), .Z(\_EXU_io_out_bits_csrOut [13] ) );
BUF_X1 \EXU/CSRControl/_3013_ ( .A(\EXU/CSRControl/csrs_4_2 [14] ), .Z(\EXU/CSRControl/_0233_ ) );
BUF_X1 \EXU/CSRControl/_3014_ ( .A(\EXU/CSRControl/csrs_3_2 [14] ), .Z(\EXU/CSRControl/_0201_ ) );
BUF_X1 \EXU/CSRControl/_3015_ ( .A(\EXU/CSRControl/csrs_2_2 [14] ), .Z(\EXU/CSRControl/_0169_ ) );
BUF_X1 \EXU/CSRControl/_3016_ ( .A(\EXU/CSRControl/csrs_0_2 [14] ), .Z(\EXU/CSRControl/_0137_ ) );
BUF_X1 \EXU/CSRControl/_3017_ ( .A(\EXU/CSRControl/_0312_ ), .Z(\_EXU_io_out_bits_csrOut [14] ) );
BUF_X1 \EXU/CSRControl/_3018_ ( .A(\EXU/CSRControl/csrs_4_2 [15] ), .Z(\EXU/CSRControl/_0234_ ) );
BUF_X1 \EXU/CSRControl/_3019_ ( .A(\EXU/CSRControl/csrs_3_2 [15] ), .Z(\EXU/CSRControl/_0202_ ) );
BUF_X1 \EXU/CSRControl/_3020_ ( .A(\EXU/CSRControl/csrs_2_2 [15] ), .Z(\EXU/CSRControl/_0170_ ) );
BUF_X1 \EXU/CSRControl/_3021_ ( .A(\EXU/CSRControl/csrs_0_2 [15] ), .Z(\EXU/CSRControl/_0138_ ) );
BUF_X1 \EXU/CSRControl/_3022_ ( .A(\EXU/CSRControl/_0313_ ), .Z(\_EXU_io_out_bits_csrOut [15] ) );
BUF_X1 \EXU/CSRControl/_3023_ ( .A(\EXU/CSRControl/csrs_4_2 [16] ), .Z(\EXU/CSRControl/_0235_ ) );
BUF_X1 \EXU/CSRControl/_3024_ ( .A(\EXU/CSRControl/csrs_3_2 [16] ), .Z(\EXU/CSRControl/_0203_ ) );
BUF_X1 \EXU/CSRControl/_3025_ ( .A(\EXU/CSRControl/csrs_2_2 [16] ), .Z(\EXU/CSRControl/_0171_ ) );
BUF_X1 \EXU/CSRControl/_3026_ ( .A(\EXU/CSRControl/csrs_0_2 [16] ), .Z(\EXU/CSRControl/_0139_ ) );
BUF_X1 \EXU/CSRControl/_3027_ ( .A(\EXU/CSRControl/_0314_ ), .Z(\_EXU_io_out_bits_csrOut [16] ) );
BUF_X1 \EXU/CSRControl/_3028_ ( .A(\EXU/CSRControl/csrs_4_2 [17] ), .Z(\EXU/CSRControl/_0236_ ) );
BUF_X1 \EXU/CSRControl/_3029_ ( .A(\EXU/CSRControl/csrs_3_2 [17] ), .Z(\EXU/CSRControl/_0204_ ) );
BUF_X1 \EXU/CSRControl/_3030_ ( .A(\EXU/CSRControl/csrs_2_2 [17] ), .Z(\EXU/CSRControl/_0172_ ) );
BUF_X1 \EXU/CSRControl/_3031_ ( .A(\EXU/CSRControl/csrs_0_2 [17] ), .Z(\EXU/CSRControl/_0140_ ) );
BUF_X1 \EXU/CSRControl/_3032_ ( .A(\EXU/CSRControl/_0315_ ), .Z(\_EXU_io_out_bits_csrOut [17] ) );
BUF_X1 \EXU/CSRControl/_3033_ ( .A(\EXU/CSRControl/csrs_4_2 [18] ), .Z(\EXU/CSRControl/_0237_ ) );
BUF_X1 \EXU/CSRControl/_3034_ ( .A(\EXU/CSRControl/csrs_3_2 [18] ), .Z(\EXU/CSRControl/_0205_ ) );
BUF_X1 \EXU/CSRControl/_3035_ ( .A(\EXU/CSRControl/csrs_2_2 [18] ), .Z(\EXU/CSRControl/_0173_ ) );
BUF_X1 \EXU/CSRControl/_3036_ ( .A(\EXU/CSRControl/csrs_0_2 [18] ), .Z(\EXU/CSRControl/_0141_ ) );
BUF_X1 \EXU/CSRControl/_3037_ ( .A(\EXU/CSRControl/_0316_ ), .Z(\_EXU_io_out_bits_csrOut [18] ) );
BUF_X1 \EXU/CSRControl/_3038_ ( .A(\EXU/CSRControl/csrs_4_2 [19] ), .Z(\EXU/CSRControl/_0238_ ) );
BUF_X1 \EXU/CSRControl/_3039_ ( .A(\EXU/CSRControl/csrs_3_2 [19] ), .Z(\EXU/CSRControl/_0206_ ) );
BUF_X1 \EXU/CSRControl/_3040_ ( .A(\EXU/CSRControl/csrs_2_2 [19] ), .Z(\EXU/CSRControl/_0174_ ) );
BUF_X1 \EXU/CSRControl/_3041_ ( .A(\EXU/CSRControl/csrs_0_2 [19] ), .Z(\EXU/CSRControl/_0142_ ) );
BUF_X1 \EXU/CSRControl/_3042_ ( .A(\EXU/CSRControl/_0317_ ), .Z(\_EXU_io_out_bits_csrOut [19] ) );
BUF_X1 \EXU/CSRControl/_3043_ ( .A(\EXU/CSRControl/csrs_4_2 [20] ), .Z(\EXU/CSRControl/_0240_ ) );
BUF_X1 \EXU/CSRControl/_3044_ ( .A(\EXU/CSRControl/csrs_3_2 [20] ), .Z(\EXU/CSRControl/_0208_ ) );
BUF_X1 \EXU/CSRControl/_3045_ ( .A(\EXU/CSRControl/csrs_2_2 [20] ), .Z(\EXU/CSRControl/_0176_ ) );
BUF_X1 \EXU/CSRControl/_3046_ ( .A(\EXU/CSRControl/csrs_0_2 [20] ), .Z(\EXU/CSRControl/_0144_ ) );
BUF_X1 \EXU/CSRControl/_3047_ ( .A(\EXU/CSRControl/_0319_ ), .Z(\_EXU_io_out_bits_csrOut [20] ) );
BUF_X1 \EXU/CSRControl/_3048_ ( .A(\EXU/CSRControl/csrs_4_2 [21] ), .Z(\EXU/CSRControl/_0241_ ) );
BUF_X1 \EXU/CSRControl/_3049_ ( .A(\EXU/CSRControl/csrs_3_2 [21] ), .Z(\EXU/CSRControl/_0209_ ) );
BUF_X1 \EXU/CSRControl/_3050_ ( .A(\EXU/CSRControl/csrs_2_2 [21] ), .Z(\EXU/CSRControl/_0177_ ) );
BUF_X1 \EXU/CSRControl/_3051_ ( .A(\EXU/CSRControl/csrs_0_2 [21] ), .Z(\EXU/CSRControl/_0145_ ) );
BUF_X1 \EXU/CSRControl/_3052_ ( .A(\EXU/CSRControl/_0320_ ), .Z(\_EXU_io_out_bits_csrOut [21] ) );
BUF_X1 \EXU/CSRControl/_3053_ ( .A(\EXU/CSRControl/csrs_4_2 [22] ), .Z(\EXU/CSRControl/_0242_ ) );
BUF_X1 \EXU/CSRControl/_3054_ ( .A(\EXU/CSRControl/csrs_3_2 [22] ), .Z(\EXU/CSRControl/_0210_ ) );
BUF_X1 \EXU/CSRControl/_3055_ ( .A(\EXU/CSRControl/csrs_2_2 [22] ), .Z(\EXU/CSRControl/_0178_ ) );
BUF_X1 \EXU/CSRControl/_3056_ ( .A(\EXU/CSRControl/csrs_0_2 [22] ), .Z(\EXU/CSRControl/_0146_ ) );
BUF_X1 \EXU/CSRControl/_3057_ ( .A(\EXU/CSRControl/_0321_ ), .Z(\_EXU_io_out_bits_csrOut [22] ) );
BUF_X1 \EXU/CSRControl/_3058_ ( .A(\EXU/CSRControl/csrs_4_2 [23] ), .Z(\EXU/CSRControl/_0243_ ) );
BUF_X1 \EXU/CSRControl/_3059_ ( .A(\EXU/CSRControl/csrs_3_2 [23] ), .Z(\EXU/CSRControl/_0211_ ) );
BUF_X1 \EXU/CSRControl/_3060_ ( .A(\EXU/CSRControl/csrs_2_2 [23] ), .Z(\EXU/CSRControl/_0179_ ) );
BUF_X1 \EXU/CSRControl/_3061_ ( .A(\EXU/CSRControl/csrs_0_2 [23] ), .Z(\EXU/CSRControl/_0147_ ) );
BUF_X1 \EXU/CSRControl/_3062_ ( .A(\EXU/CSRControl/_0322_ ), .Z(\_EXU_io_out_bits_csrOut [23] ) );
BUF_X1 \EXU/CSRControl/_3063_ ( .A(\EXU/CSRControl/csrs_4_2 [24] ), .Z(\EXU/CSRControl/_0244_ ) );
BUF_X1 \EXU/CSRControl/_3064_ ( .A(\EXU/CSRControl/csrs_3_2 [24] ), .Z(\EXU/CSRControl/_0212_ ) );
BUF_X1 \EXU/CSRControl/_3065_ ( .A(\EXU/CSRControl/csrs_2_2 [24] ), .Z(\EXU/CSRControl/_0180_ ) );
BUF_X1 \EXU/CSRControl/_3066_ ( .A(\EXU/CSRControl/csrs_0_2 [24] ), .Z(\EXU/CSRControl/_0148_ ) );
BUF_X1 \EXU/CSRControl/_3067_ ( .A(\EXU/CSRControl/_0323_ ), .Z(\_EXU_io_out_bits_csrOut [24] ) );
BUF_X1 \EXU/CSRControl/_3068_ ( .A(\EXU/CSRControl/csrs_4_2 [25] ), .Z(\EXU/CSRControl/_0245_ ) );
BUF_X1 \EXU/CSRControl/_3069_ ( .A(\EXU/CSRControl/csrs_3_2 [25] ), .Z(\EXU/CSRControl/_0213_ ) );
BUF_X1 \EXU/CSRControl/_3070_ ( .A(\EXU/CSRControl/csrs_2_2 [25] ), .Z(\EXU/CSRControl/_0181_ ) );
BUF_X1 \EXU/CSRControl/_3071_ ( .A(\EXU/CSRControl/csrs_0_2 [25] ), .Z(\EXU/CSRControl/_0149_ ) );
BUF_X1 \EXU/CSRControl/_3072_ ( .A(\EXU/CSRControl/_0324_ ), .Z(\_EXU_io_out_bits_csrOut [25] ) );
BUF_X1 \EXU/CSRControl/_3073_ ( .A(\EXU/CSRControl/csrs_4_2 [26] ), .Z(\EXU/CSRControl/_0246_ ) );
BUF_X1 \EXU/CSRControl/_3074_ ( .A(\EXU/CSRControl/csrs_3_2 [26] ), .Z(\EXU/CSRControl/_0214_ ) );
BUF_X1 \EXU/CSRControl/_3075_ ( .A(\EXU/CSRControl/csrs_2_2 [26] ), .Z(\EXU/CSRControl/_0182_ ) );
BUF_X1 \EXU/CSRControl/_3076_ ( .A(\EXU/CSRControl/csrs_0_2 [26] ), .Z(\EXU/CSRControl/_0150_ ) );
BUF_X1 \EXU/CSRControl/_3077_ ( .A(\EXU/CSRControl/_0325_ ), .Z(\_EXU_io_out_bits_csrOut [26] ) );
BUF_X1 \EXU/CSRControl/_3078_ ( .A(\EXU/CSRControl/csrs_4_2 [27] ), .Z(\EXU/CSRControl/_0247_ ) );
BUF_X1 \EXU/CSRControl/_3079_ ( .A(\EXU/CSRControl/csrs_3_2 [27] ), .Z(\EXU/CSRControl/_0215_ ) );
BUF_X1 \EXU/CSRControl/_3080_ ( .A(\EXU/CSRControl/csrs_2_2 [27] ), .Z(\EXU/CSRControl/_0183_ ) );
BUF_X1 \EXU/CSRControl/_3081_ ( .A(\EXU/CSRControl/csrs_0_2 [27] ), .Z(\EXU/CSRControl/_0151_ ) );
BUF_X1 \EXU/CSRControl/_3082_ ( .A(\EXU/CSRControl/_0326_ ), .Z(\_EXU_io_out_bits_csrOut [27] ) );
BUF_X1 \EXU/CSRControl/_3083_ ( .A(\EXU/CSRControl/csrs_4_2 [28] ), .Z(\EXU/CSRControl/_0248_ ) );
BUF_X1 \EXU/CSRControl/_3084_ ( .A(\EXU/CSRControl/csrs_3_2 [28] ), .Z(\EXU/CSRControl/_0216_ ) );
BUF_X1 \EXU/CSRControl/_3085_ ( .A(\EXU/CSRControl/csrs_2_2 [28] ), .Z(\EXU/CSRControl/_0184_ ) );
BUF_X1 \EXU/CSRControl/_3086_ ( .A(\EXU/CSRControl/csrs_0_2 [28] ), .Z(\EXU/CSRControl/_0152_ ) );
BUF_X1 \EXU/CSRControl/_3087_ ( .A(\EXU/CSRControl/_0327_ ), .Z(\_EXU_io_out_bits_csrOut [28] ) );
BUF_X1 \EXU/CSRControl/_3088_ ( .A(\EXU/CSRControl/csrs_4_2 [29] ), .Z(\EXU/CSRControl/_0249_ ) );
BUF_X1 \EXU/CSRControl/_3089_ ( .A(\EXU/CSRControl/csrs_3_2 [29] ), .Z(\EXU/CSRControl/_0217_ ) );
BUF_X1 \EXU/CSRControl/_3090_ ( .A(\EXU/CSRControl/csrs_2_2 [29] ), .Z(\EXU/CSRControl/_0185_ ) );
BUF_X1 \EXU/CSRControl/_3091_ ( .A(\EXU/CSRControl/csrs_0_2 [29] ), .Z(\EXU/CSRControl/_0153_ ) );
BUF_X1 \EXU/CSRControl/_3092_ ( .A(\EXU/CSRControl/_0328_ ), .Z(\_EXU_io_out_bits_csrOut [29] ) );
BUF_X1 \EXU/CSRControl/_3093_ ( .A(\EXU/CSRControl/csrs_4_2 [30] ), .Z(\EXU/CSRControl/_0251_ ) );
BUF_X1 \EXU/CSRControl/_3094_ ( .A(\EXU/CSRControl/csrs_3_2 [30] ), .Z(\EXU/CSRControl/_0219_ ) );
BUF_X1 \EXU/CSRControl/_3095_ ( .A(\EXU/CSRControl/csrs_2_2 [30] ), .Z(\EXU/CSRControl/_0187_ ) );
BUF_X1 \EXU/CSRControl/_3096_ ( .A(\EXU/CSRControl/csrs_0_2 [30] ), .Z(\EXU/CSRControl/_0155_ ) );
BUF_X1 \EXU/CSRControl/_3097_ ( .A(\EXU/CSRControl/_0330_ ), .Z(\_EXU_io_out_bits_csrOut [30] ) );
BUF_X1 \EXU/CSRControl/_3098_ ( .A(\EXU/CSRControl/csrs_4_2 [31] ), .Z(\EXU/CSRControl/_0252_ ) );
BUF_X1 \EXU/CSRControl/_3099_ ( .A(\EXU/CSRControl/csrs_3_2 [31] ), .Z(\EXU/CSRControl/_0220_ ) );
BUF_X1 \EXU/CSRControl/_3100_ ( .A(\EXU/CSRControl/csrs_2_2 [31] ), .Z(\EXU/CSRControl/_0188_ ) );
BUF_X1 \EXU/CSRControl/_3101_ ( .A(\EXU/CSRControl/csrs_0_2 [31] ), .Z(\EXU/CSRControl/_0156_ ) );
BUF_X1 \EXU/CSRControl/_3102_ ( .A(\EXU/CSRControl/_0331_ ), .Z(\_EXU_io_out_bits_csrOut [31] ) );
BUF_X1 \EXU/CSRControl/_3103_ ( .A(\EXU/_0035_ ), .Z(\EXU/CSRControl/_0275_ ) );
BUF_X1 \EXU/CSRControl/_3104_ ( .A(\EXU/_0046_ ), .Z(\EXU/CSRControl/_0286_ ) );
BUF_X1 \EXU/CSRControl/_3105_ ( .A(\EXU/_0057_ ), .Z(\EXU/CSRControl/_0297_ ) );
BUF_X1 \EXU/CSRControl/_3106_ ( .A(\EXU/_0060_ ), .Z(\EXU/CSRControl/_0300_ ) );
BUF_X1 \EXU/CSRControl/_3107_ ( .A(\EXU/_0061_ ), .Z(\EXU/CSRControl/_0301_ ) );
BUF_X1 \EXU/CSRControl/_3108_ ( .A(\EXU/_0062_ ), .Z(\EXU/CSRControl/_0302_ ) );
BUF_X1 \EXU/CSRControl/_3109_ ( .A(\EXU/_0063_ ), .Z(\EXU/CSRControl/_0303_ ) );
BUF_X1 \EXU/CSRControl/_3110_ ( .A(\EXU/_0064_ ), .Z(\EXU/CSRControl/_0304_ ) );
BUF_X1 \EXU/CSRControl/_3111_ ( .A(\EXU/_0065_ ), .Z(\EXU/CSRControl/_0305_ ) );
BUF_X1 \EXU/CSRControl/_3112_ ( .A(\EXU/_0066_ ), .Z(\EXU/CSRControl/_0306_ ) );
BUF_X1 \EXU/CSRControl/_3113_ ( .A(\EXU/_0036_ ), .Z(\EXU/CSRControl/_0276_ ) );
BUF_X1 \EXU/CSRControl/_3114_ ( .A(\EXU/_0037_ ), .Z(\EXU/CSRControl/_0277_ ) );
BUF_X1 \EXU/CSRControl/_3115_ ( .A(\EXU/_0038_ ), .Z(\EXU/CSRControl/_0278_ ) );
BUF_X1 \EXU/CSRControl/_3116_ ( .A(\EXU/_0039_ ), .Z(\EXU/CSRControl/_0279_ ) );
BUF_X1 \EXU/CSRControl/_3117_ ( .A(\EXU/_0040_ ), .Z(\EXU/CSRControl/_0280_ ) );
BUF_X1 \EXU/CSRControl/_3118_ ( .A(\EXU/_0041_ ), .Z(\EXU/CSRControl/_0281_ ) );
BUF_X1 \EXU/CSRControl/_3119_ ( .A(\EXU/_0042_ ), .Z(\EXU/CSRControl/_0282_ ) );
BUF_X1 \EXU/CSRControl/_3120_ ( .A(\EXU/_0043_ ), .Z(\EXU/CSRControl/_0283_ ) );
BUF_X1 \EXU/CSRControl/_3121_ ( .A(\EXU/_0044_ ), .Z(\EXU/CSRControl/_0284_ ) );
BUF_X1 \EXU/CSRControl/_3122_ ( .A(\EXU/_0045_ ), .Z(\EXU/CSRControl/_0285_ ) );
BUF_X1 \EXU/CSRControl/_3123_ ( .A(\EXU/_0047_ ), .Z(\EXU/CSRControl/_0287_ ) );
BUF_X1 \EXU/CSRControl/_3124_ ( .A(\EXU/_0048_ ), .Z(\EXU/CSRControl/_0288_ ) );
BUF_X1 \EXU/CSRControl/_3125_ ( .A(\EXU/_0049_ ), .Z(\EXU/CSRControl/_0289_ ) );
BUF_X1 \EXU/CSRControl/_3126_ ( .A(\EXU/_0050_ ), .Z(\EXU/CSRControl/_0290_ ) );
BUF_X1 \EXU/CSRControl/_3127_ ( .A(\EXU/_0051_ ), .Z(\EXU/CSRControl/_0291_ ) );
BUF_X1 \EXU/CSRControl/_3128_ ( .A(\EXU/_0052_ ), .Z(\EXU/CSRControl/_0292_ ) );
BUF_X1 \EXU/CSRControl/_3129_ ( .A(\EXU/_0053_ ), .Z(\EXU/CSRControl/_0293_ ) );
BUF_X1 \EXU/CSRControl/_3130_ ( .A(\EXU/_0054_ ), .Z(\EXU/CSRControl/_0294_ ) );
BUF_X1 \EXU/CSRControl/_3131_ ( .A(\EXU/_0055_ ), .Z(\EXU/CSRControl/_0295_ ) );
BUF_X1 \EXU/CSRControl/_3132_ ( .A(\EXU/_0056_ ), .Z(\EXU/CSRControl/_0296_ ) );
BUF_X1 \EXU/CSRControl/_3133_ ( .A(\EXU/_0058_ ), .Z(\EXU/CSRControl/_0298_ ) );
BUF_X1 \EXU/CSRControl/_3134_ ( .A(\EXU/_0059_ ), .Z(\EXU/CSRControl/_0299_ ) );
BUF_X1 \EXU/CSRControl/_3135_ ( .A(\EXU/CSRControl/priv [0] ), .Z(\EXU/CSRControl/_1372_ ) );
BUF_X1 \EXU/CSRControl/_3136_ ( .A(\EXU/CSRControl/priv [1] ), .Z(\EXU/CSRControl/_1373_ ) );
BUF_X1 \EXU/CSRControl/_3137_ ( .A(\EXU/in_pc [0] ), .Z(\EXU/CSRControl/_0339_ ) );
BUF_X1 \EXU/CSRControl/_3138_ ( .A(\EXU/in_pc [1] ), .Z(\EXU/CSRControl/_0350_ ) );
BUF_X1 \EXU/CSRControl/_3139_ ( .A(\EXU/in_pc [2] ), .Z(\EXU/CSRControl/_0361_ ) );
BUF_X1 \EXU/CSRControl/_3140_ ( .A(\EXU/in_pc [3] ), .Z(\EXU/CSRControl/_0364_ ) );
BUF_X1 \EXU/CSRControl/_3141_ ( .A(\EXU/in_pc [4] ), .Z(\EXU/CSRControl/_0365_ ) );
BUF_X1 \EXU/CSRControl/_3142_ ( .A(\EXU/in_pc [5] ), .Z(\EXU/CSRControl/_0366_ ) );
BUF_X1 \EXU/CSRControl/_3143_ ( .A(\EXU/in_pc [6] ), .Z(\EXU/CSRControl/_0367_ ) );
BUF_X1 \EXU/CSRControl/_3144_ ( .A(\EXU/in_pc [7] ), .Z(\EXU/CSRControl/_0368_ ) );
BUF_X1 \EXU/CSRControl/_3145_ ( .A(\EXU/in_pc [8] ), .Z(\EXU/CSRControl/_0369_ ) );
BUF_X1 \EXU/CSRControl/_3146_ ( .A(\EXU/in_pc [9] ), .Z(\EXU/CSRControl/_0370_ ) );
BUF_X1 \EXU/CSRControl/_3147_ ( .A(\EXU/in_pc [10] ), .Z(\EXU/CSRControl/_0340_ ) );
BUF_X1 \EXU/CSRControl/_3148_ ( .A(\EXU/in_pc [11] ), .Z(\EXU/CSRControl/_0341_ ) );
BUF_X1 \EXU/CSRControl/_3149_ ( .A(\EXU/in_pc [12] ), .Z(\EXU/CSRControl/_0342_ ) );
BUF_X1 \EXU/CSRControl/_3150_ ( .A(\EXU/in_pc [13] ), .Z(\EXU/CSRControl/_0343_ ) );
BUF_X1 \EXU/CSRControl/_3151_ ( .A(\EXU/in_pc [14] ), .Z(\EXU/CSRControl/_0344_ ) );
BUF_X1 \EXU/CSRControl/_3152_ ( .A(\EXU/in_pc [15] ), .Z(\EXU/CSRControl/_0345_ ) );
BUF_X1 \EXU/CSRControl/_3153_ ( .A(\EXU/in_pc [16] ), .Z(\EXU/CSRControl/_0346_ ) );
BUF_X1 \EXU/CSRControl/_3154_ ( .A(\EXU/in_pc [17] ), .Z(\EXU/CSRControl/_0347_ ) );
BUF_X1 \EXU/CSRControl/_3155_ ( .A(\EXU/in_pc [18] ), .Z(\EXU/CSRControl/_0348_ ) );
BUF_X1 \EXU/CSRControl/_3156_ ( .A(\EXU/in_pc [19] ), .Z(\EXU/CSRControl/_0349_ ) );
BUF_X1 \EXU/CSRControl/_3157_ ( .A(\EXU/in_pc [20] ), .Z(\EXU/CSRControl/_0351_ ) );
BUF_X1 \EXU/CSRControl/_3158_ ( .A(\EXU/in_pc [21] ), .Z(\EXU/CSRControl/_0352_ ) );
BUF_X1 \EXU/CSRControl/_3159_ ( .A(\EXU/in_pc [22] ), .Z(\EXU/CSRControl/_0353_ ) );
BUF_X1 \EXU/CSRControl/_3160_ ( .A(\EXU/in_pc [23] ), .Z(\EXU/CSRControl/_0354_ ) );
BUF_X1 \EXU/CSRControl/_3161_ ( .A(\EXU/in_pc [24] ), .Z(\EXU/CSRControl/_0355_ ) );
BUF_X1 \EXU/CSRControl/_3162_ ( .A(\EXU/in_pc [25] ), .Z(\EXU/CSRControl/_0356_ ) );
BUF_X1 \EXU/CSRControl/_3163_ ( .A(\EXU/in_pc [26] ), .Z(\EXU/CSRControl/_0357_ ) );
BUF_X1 \EXU/CSRControl/_3164_ ( .A(\EXU/in_pc [27] ), .Z(\EXU/CSRControl/_0358_ ) );
BUF_X1 \EXU/CSRControl/_3165_ ( .A(\EXU/in_pc [28] ), .Z(\EXU/CSRControl/_0359_ ) );
BUF_X1 \EXU/CSRControl/_3166_ ( .A(\EXU/in_pc [29] ), .Z(\EXU/CSRControl/_0360_ ) );
BUF_X1 \EXU/CSRControl/_3167_ ( .A(\EXU/in_pc [30] ), .Z(\EXU/CSRControl/_0362_ ) );
BUF_X1 \EXU/CSRControl/_3168_ ( .A(\EXU/in_pc [31] ), .Z(\EXU/CSRControl/_0363_ ) );
BUF_X1 \EXU/CSRControl/_3169_ ( .A(\EXU/CSRControl/_0000_ ), .Z(\EXU/CSRControl/_0001_ ) );
BUF_X1 \EXU/CSRControl/_3170_ ( .A(\EXU/CSRControl/_0002_ ), .Z(\EXU/CSRControl/_1504_ ) );
BUF_X1 \EXU/CSRControl/_3171_ ( .A(\EXU/CSRControl/_0003_ ), .Z(\EXU/CSRControl/_1505_ ) );
BUF_X1 \EXU/CSRControl/_3172_ ( .A(\EXU/CSRControl/_0004_ ), .Z(\EXU/CSRControl/_1506_ ) );
BUF_X1 \EXU/CSRControl/_3173_ ( .A(\EXU/CSRControl/_0005_ ), .Z(\EXU/CSRControl/_1507_ ) );
BUF_X1 \EXU/CSRControl/_3174_ ( .A(\EXU/CSRControl/_0006_ ), .Z(\EXU/CSRControl/_1508_ ) );
BUF_X1 \EXU/CSRControl/_3175_ ( .A(\EXU/CSRControl/_0007_ ), .Z(\EXU/CSRControl/_1509_ ) );
BUF_X1 \EXU/CSRControl/_3176_ ( .A(\EXU/CSRControl/_0008_ ), .Z(\EXU/CSRControl/_1510_ ) );
BUF_X1 \EXU/CSRControl/_3177_ ( .A(\EXU/CSRControl/_0009_ ), .Z(\EXU/CSRControl/_1511_ ) );
BUF_X1 \EXU/CSRControl/_3178_ ( .A(\EXU/CSRControl/_0010_ ), .Z(\EXU/CSRControl/_1512_ ) );
BUF_X1 \EXU/CSRControl/_3179_ ( .A(\EXU/CSRControl/_0011_ ), .Z(\EXU/CSRControl/_1513_ ) );
BUF_X1 \EXU/CSRControl/_3180_ ( .A(\EXU/CSRControl/_0012_ ), .Z(\EXU/CSRControl/_1514_ ) );
BUF_X1 \EXU/CSRControl/_3181_ ( .A(\EXU/CSRControl/_0013_ ), .Z(\EXU/CSRControl/_1515_ ) );
BUF_X1 \EXU/CSRControl/_3182_ ( .A(\EXU/CSRControl/_0014_ ), .Z(\EXU/CSRControl/_1516_ ) );
BUF_X1 \EXU/CSRControl/_3183_ ( .A(\EXU/CSRControl/_0015_ ), .Z(\EXU/CSRControl/_1517_ ) );
BUF_X1 \EXU/CSRControl/_3184_ ( .A(\EXU/CSRControl/_0016_ ), .Z(\EXU/CSRControl/_1518_ ) );
BUF_X1 \EXU/CSRControl/_3185_ ( .A(\EXU/CSRControl/_0017_ ), .Z(\EXU/CSRControl/_1519_ ) );
BUF_X1 \EXU/CSRControl/_3186_ ( .A(\EXU/CSRControl/_0018_ ), .Z(\EXU/CSRControl/_1520_ ) );
BUF_X1 \EXU/CSRControl/_3187_ ( .A(\EXU/CSRControl/_0019_ ), .Z(\EXU/CSRControl/_1521_ ) );
BUF_X1 \EXU/CSRControl/_3188_ ( .A(\EXU/CSRControl/_0020_ ), .Z(\EXU/CSRControl/_1522_ ) );
BUF_X1 \EXU/CSRControl/_3189_ ( .A(\EXU/CSRControl/_0021_ ), .Z(\EXU/CSRControl/_1523_ ) );
BUF_X1 \EXU/CSRControl/_3190_ ( .A(\EXU/CSRControl/_0022_ ), .Z(\EXU/CSRControl/_1524_ ) );
BUF_X1 \EXU/CSRControl/_3191_ ( .A(\EXU/CSRControl/_0023_ ), .Z(\EXU/CSRControl/_1525_ ) );
BUF_X1 \EXU/CSRControl/_3192_ ( .A(\EXU/CSRControl/_0024_ ), .Z(\EXU/CSRControl/_1526_ ) );
BUF_X1 \EXU/CSRControl/_3193_ ( .A(\EXU/CSRControl/_0025_ ), .Z(\EXU/CSRControl/_1527_ ) );
BUF_X1 \EXU/CSRControl/_3194_ ( .A(\EXU/CSRControl/_0026_ ), .Z(\EXU/CSRControl/_1528_ ) );
BUF_X1 \EXU/CSRControl/_3195_ ( .A(\EXU/CSRControl/_0027_ ), .Z(\EXU/CSRControl/_1529_ ) );
BUF_X1 \EXU/CSRControl/_3196_ ( .A(\EXU/CSRControl/_0028_ ), .Z(\EXU/CSRControl/_1530_ ) );
BUF_X1 \EXU/CSRControl/_3197_ ( .A(\EXU/CSRControl/_0029_ ), .Z(\EXU/CSRControl/_1531_ ) );
BUF_X1 \EXU/CSRControl/_3198_ ( .A(\EXU/CSRControl/_0030_ ), .Z(\EXU/CSRControl/_1532_ ) );
BUF_X1 \EXU/CSRControl/_3199_ ( .A(\EXU/CSRControl/_0031_ ), .Z(\EXU/CSRControl/_1533_ ) );
BUF_X1 \EXU/CSRControl/_3200_ ( .A(\EXU/CSRControl/_0032_ ), .Z(\EXU/CSRControl/_1534_ ) );
BUF_X1 \EXU/CSRControl/_3201_ ( .A(\EXU/CSRControl/_0033_ ), .Z(\EXU/CSRControl/_1535_ ) );
BUF_X1 \EXU/CSRControl/_3202_ ( .A(\EXU/CSRControl/_0034_ ), .Z(\EXU/CSRControl/_1536_ ) );
BUF_X1 \EXU/CSRControl/_3203_ ( .A(\EXU/CSRControl/_0035_ ), .Z(\EXU/CSRControl/_1537_ ) );
BUF_X1 \EXU/CSRControl/_3204_ ( .A(\EXU/CSRControl/_0036_ ), .Z(\EXU/CSRControl/_1538_ ) );
BUF_X1 \EXU/CSRControl/_3205_ ( .A(\EXU/CSRControl/_0037_ ), .Z(\EXU/CSRControl/_1539_ ) );
BUF_X1 \EXU/CSRControl/_3206_ ( .A(\EXU/CSRControl/_0038_ ), .Z(\EXU/CSRControl/_1540_ ) );
BUF_X1 \EXU/CSRControl/_3207_ ( .A(\EXU/CSRControl/_0039_ ), .Z(\EXU/CSRControl/_1541_ ) );
BUF_X1 \EXU/CSRControl/_3208_ ( .A(\EXU/CSRControl/_0040_ ), .Z(\EXU/CSRControl/_1542_ ) );
BUF_X1 \EXU/CSRControl/_3209_ ( .A(\EXU/CSRControl/_0041_ ), .Z(\EXU/CSRControl/_1543_ ) );
BUF_X1 \EXU/CSRControl/_3210_ ( .A(\EXU/CSRControl/_0042_ ), .Z(\EXU/CSRControl/_1544_ ) );
BUF_X1 \EXU/CSRControl/_3211_ ( .A(\EXU/CSRControl/_0043_ ), .Z(\EXU/CSRControl/_1545_ ) );
BUF_X1 \EXU/CSRControl/_3212_ ( .A(\EXU/CSRControl/_0044_ ), .Z(\EXU/CSRControl/_1546_ ) );
BUF_X1 \EXU/CSRControl/_3213_ ( .A(\EXU/CSRControl/_0045_ ), .Z(\EXU/CSRControl/_1547_ ) );
BUF_X1 \EXU/CSRControl/_3214_ ( .A(\EXU/CSRControl/_0046_ ), .Z(\EXU/CSRControl/_1548_ ) );
BUF_X1 \EXU/CSRControl/_3215_ ( .A(\EXU/CSRControl/_0047_ ), .Z(\EXU/CSRControl/_1549_ ) );
BUF_X1 \EXU/CSRControl/_3216_ ( .A(\EXU/CSRControl/_0048_ ), .Z(\EXU/CSRControl/_1550_ ) );
BUF_X1 \EXU/CSRControl/_3217_ ( .A(\EXU/CSRControl/_0049_ ), .Z(\EXU/CSRControl/_1551_ ) );
BUF_X1 \EXU/CSRControl/_3218_ ( .A(\EXU/CSRControl/_0050_ ), .Z(\EXU/CSRControl/_1552_ ) );
BUF_X1 \EXU/CSRControl/_3219_ ( .A(\EXU/CSRControl/_0051_ ), .Z(\EXU/CSRControl/_1553_ ) );
BUF_X1 \EXU/CSRControl/_3220_ ( .A(\EXU/CSRControl/_0052_ ), .Z(\EXU/CSRControl/_1554_ ) );
BUF_X1 \EXU/CSRControl/_3221_ ( .A(\EXU/CSRControl/_0053_ ), .Z(\EXU/CSRControl/_1555_ ) );
BUF_X1 \EXU/CSRControl/_3222_ ( .A(\EXU/CSRControl/_0054_ ), .Z(\EXU/CSRControl/_1556_ ) );
BUF_X1 \EXU/CSRControl/_3223_ ( .A(\EXU/CSRControl/_0055_ ), .Z(\EXU/CSRControl/_1557_ ) );
BUF_X1 \EXU/CSRControl/_3224_ ( .A(\EXU/CSRControl/_0056_ ), .Z(\EXU/CSRControl/_1558_ ) );
BUF_X1 \EXU/CSRControl/_3225_ ( .A(\EXU/CSRControl/_0057_ ), .Z(\EXU/CSRControl/_1559_ ) );
BUF_X1 \EXU/CSRControl/_3226_ ( .A(\EXU/CSRControl/_0058_ ), .Z(\EXU/CSRControl/_1560_ ) );
BUF_X1 \EXU/CSRControl/_3227_ ( .A(\EXU/CSRControl/_0059_ ), .Z(\EXU/CSRControl/_1561_ ) );
BUF_X1 \EXU/CSRControl/_3228_ ( .A(\EXU/CSRControl/_0060_ ), .Z(\EXU/CSRControl/_1562_ ) );
BUF_X1 \EXU/CSRControl/_3229_ ( .A(\EXU/CSRControl/_0061_ ), .Z(\EXU/CSRControl/_1563_ ) );
BUF_X1 \EXU/CSRControl/_3230_ ( .A(\EXU/CSRControl/_0062_ ), .Z(\EXU/CSRControl/_1564_ ) );
BUF_X1 \EXU/CSRControl/_3231_ ( .A(\EXU/CSRControl/_0063_ ), .Z(\EXU/CSRControl/_1565_ ) );
BUF_X1 \EXU/CSRControl/_3232_ ( .A(\EXU/CSRControl/_0064_ ), .Z(\EXU/CSRControl/_1566_ ) );
BUF_X1 \EXU/CSRControl/_3233_ ( .A(\EXU/CSRControl/_0065_ ), .Z(\EXU/CSRControl/_1567_ ) );
BUF_X1 \EXU/CSRControl/_3234_ ( .A(\EXU/CSRControl/_0066_ ), .Z(\EXU/CSRControl/_1568_ ) );
BUF_X1 \EXU/CSRControl/_3235_ ( .A(\EXU/CSRControl/_0067_ ), .Z(\EXU/CSRControl/_1569_ ) );
BUF_X1 \EXU/CSRControl/_3236_ ( .A(\EXU/CSRControl/_0068_ ), .Z(\EXU/CSRControl/_1570_ ) );
BUF_X1 \EXU/CSRControl/_3237_ ( .A(\EXU/CSRControl/_0069_ ), .Z(\EXU/CSRControl/_1571_ ) );
BUF_X1 \EXU/CSRControl/_3238_ ( .A(\EXU/CSRControl/_0070_ ), .Z(\EXU/CSRControl/_1572_ ) );
BUF_X1 \EXU/CSRControl/_3239_ ( .A(\EXU/CSRControl/_0071_ ), .Z(\EXU/CSRControl/_1573_ ) );
BUF_X1 \EXU/CSRControl/_3240_ ( .A(\EXU/CSRControl/_0072_ ), .Z(\EXU/CSRControl/_1574_ ) );
BUF_X1 \EXU/CSRControl/_3241_ ( .A(\EXU/CSRControl/_0073_ ), .Z(\EXU/CSRControl/_1575_ ) );
BUF_X1 \EXU/CSRControl/_3242_ ( .A(\EXU/CSRControl/_0074_ ), .Z(\EXU/CSRControl/_1576_ ) );
BUF_X1 \EXU/CSRControl/_3243_ ( .A(\EXU/CSRControl/_0075_ ), .Z(\EXU/CSRControl/_1577_ ) );
BUF_X1 \EXU/CSRControl/_3244_ ( .A(\EXU/CSRControl/_0076_ ), .Z(\EXU/CSRControl/_1578_ ) );
BUF_X1 \EXU/CSRControl/_3245_ ( .A(\EXU/CSRControl/_0077_ ), .Z(\EXU/CSRControl/_1579_ ) );
BUF_X1 \EXU/CSRControl/_3246_ ( .A(\EXU/CSRControl/_0078_ ), .Z(\EXU/CSRControl/_1580_ ) );
BUF_X1 \EXU/CSRControl/_3247_ ( .A(\EXU/CSRControl/_0079_ ), .Z(\EXU/CSRControl/_1581_ ) );
BUF_X1 \EXU/CSRControl/_3248_ ( .A(\EXU/CSRControl/_0080_ ), .Z(\EXU/CSRControl/_1582_ ) );
BUF_X1 \EXU/CSRControl/_3249_ ( .A(\EXU/CSRControl/_0081_ ), .Z(\EXU/CSRControl/_1583_ ) );
BUF_X1 \EXU/CSRControl/_3250_ ( .A(\EXU/CSRControl/_0082_ ), .Z(\EXU/CSRControl/_1584_ ) );
BUF_X1 \EXU/CSRControl/_3251_ ( .A(\EXU/CSRControl/_0083_ ), .Z(\EXU/CSRControl/_1585_ ) );
BUF_X1 \EXU/CSRControl/_3252_ ( .A(\EXU/CSRControl/_0084_ ), .Z(\EXU/CSRControl/_1586_ ) );
BUF_X1 \EXU/CSRControl/_3253_ ( .A(\EXU/CSRControl/_0085_ ), .Z(\EXU/CSRControl/_1587_ ) );
BUF_X1 \EXU/CSRControl/_3254_ ( .A(\EXU/CSRControl/_0086_ ), .Z(\EXU/CSRControl/_1588_ ) );
BUF_X1 \EXU/CSRControl/_3255_ ( .A(\EXU/CSRControl/_0087_ ), .Z(\EXU/CSRControl/_1589_ ) );
BUF_X1 \EXU/CSRControl/_3256_ ( .A(\EXU/CSRControl/_0088_ ), .Z(\EXU/CSRControl/_1590_ ) );
BUF_X1 \EXU/CSRControl/_3257_ ( .A(\EXU/CSRControl/_0089_ ), .Z(\EXU/CSRControl/_1591_ ) );
BUF_X1 \EXU/CSRControl/_3258_ ( .A(\EXU/CSRControl/_0090_ ), .Z(\EXU/CSRControl/_1592_ ) );
BUF_X1 \EXU/CSRControl/_3259_ ( .A(\EXU/CSRControl/_0091_ ), .Z(\EXU/CSRControl/_1593_ ) );
BUF_X1 \EXU/CSRControl/_3260_ ( .A(\EXU/CSRControl/_0092_ ), .Z(\EXU/CSRControl/_1594_ ) );
BUF_X1 \EXU/CSRControl/_3261_ ( .A(\EXU/CSRControl/_0093_ ), .Z(\EXU/CSRControl/_1595_ ) );
BUF_X1 \EXU/CSRControl/_3262_ ( .A(\EXU/CSRControl/_0094_ ), .Z(\EXU/CSRControl/_1596_ ) );
BUF_X1 \EXU/CSRControl/_3263_ ( .A(\EXU/CSRControl/_0095_ ), .Z(\EXU/CSRControl/_1597_ ) );
BUF_X1 \EXU/CSRControl/_3264_ ( .A(\EXU/CSRControl/_0096_ ), .Z(\EXU/CSRControl/_1598_ ) );
BUF_X1 \EXU/CSRControl/_3265_ ( .A(\EXU/CSRControl/_0097_ ), .Z(\EXU/CSRControl/_1599_ ) );
BUF_X1 \EXU/CSRControl/_3266_ ( .A(\EXU/CSRControl/_0098_ ), .Z(\EXU/CSRControl/_1600_ ) );
BUF_X1 \EXU/CSRControl/_3267_ ( .A(\EXU/CSRControl/_0099_ ), .Z(\EXU/CSRControl/_1601_ ) );
BUF_X1 \EXU/CSRControl/_3268_ ( .A(\EXU/CSRControl/_0100_ ), .Z(\EXU/CSRControl/_1602_ ) );
BUF_X1 \EXU/CSRControl/_3269_ ( .A(\EXU/CSRControl/_0101_ ), .Z(\EXU/CSRControl/_1603_ ) );
BUF_X1 \EXU/CSRControl/_3270_ ( .A(\EXU/CSRControl/_0102_ ), .Z(\EXU/CSRControl/_1604_ ) );
BUF_X1 \EXU/CSRControl/_3271_ ( .A(\EXU/CSRControl/_0103_ ), .Z(\EXU/CSRControl/_1605_ ) );
BUF_X1 \EXU/CSRControl/_3272_ ( .A(\EXU/CSRControl/_0104_ ), .Z(\EXU/CSRControl/_1606_ ) );
BUF_X1 \EXU/CSRControl/_3273_ ( .A(\EXU/CSRControl/_0105_ ), .Z(\EXU/CSRControl/_1607_ ) );
BUF_X1 \EXU/CSRControl/_3274_ ( .A(\EXU/CSRControl/_0106_ ), .Z(\EXU/CSRControl/_1608_ ) );
BUF_X1 \EXU/CSRControl/_3275_ ( .A(\EXU/CSRControl/_0107_ ), .Z(\EXU/CSRControl/_1609_ ) );
BUF_X1 \EXU/CSRControl/_3276_ ( .A(\EXU/CSRControl/_0108_ ), .Z(\EXU/CSRControl/_1610_ ) );
BUF_X1 \EXU/CSRControl/_3277_ ( .A(\EXU/CSRControl/_0109_ ), .Z(\EXU/CSRControl/_1611_ ) );
BUF_X1 \EXU/CSRControl/_3278_ ( .A(\EXU/CSRControl/_0110_ ), .Z(\EXU/CSRControl/_1612_ ) );
BUF_X1 \EXU/CSRControl/_3279_ ( .A(\EXU/CSRControl/_0111_ ), .Z(\EXU/CSRControl/_1613_ ) );
BUF_X1 \EXU/CSRControl/_3280_ ( .A(\EXU/CSRControl/_0112_ ), .Z(\EXU/CSRControl/_1614_ ) );
BUF_X1 \EXU/CSRControl/_3281_ ( .A(\EXU/CSRControl/_0113_ ), .Z(\EXU/CSRControl/_1615_ ) );
BUF_X1 \EXU/CSRControl/_3282_ ( .A(\EXU/CSRControl/_0114_ ), .Z(\EXU/CSRControl/_1616_ ) );
BUF_X1 \EXU/CSRControl/_3283_ ( .A(\EXU/CSRControl/_0115_ ), .Z(\EXU/CSRControl/_1617_ ) );
BUF_X1 \EXU/CSRControl/_3284_ ( .A(\EXU/CSRControl/_0116_ ), .Z(\EXU/CSRControl/_1618_ ) );
BUF_X1 \EXU/CSRControl/_3285_ ( .A(\EXU/CSRControl/_0117_ ), .Z(\EXU/CSRControl/_1619_ ) );
BUF_X1 \EXU/CSRControl/_3286_ ( .A(\EXU/CSRControl/_0118_ ), .Z(\EXU/CSRControl/_1620_ ) );
BUF_X1 \EXU/CSRControl/_3287_ ( .A(\EXU/CSRControl/_0119_ ), .Z(\EXU/CSRControl/_1621_ ) );
BUF_X1 \EXU/CSRControl/_3288_ ( .A(\EXU/CSRControl/_0120_ ), .Z(\EXU/CSRControl/_1622_ ) );
BUF_X1 \EXU/CSRControl/_3289_ ( .A(\EXU/CSRControl/_0121_ ), .Z(\EXU/CSRControl/_1623_ ) );
BUF_X1 \EXU/CSRControl/_3290_ ( .A(\EXU/CSRControl/_0122_ ), .Z(\EXU/CSRControl/_1624_ ) );
BUF_X1 \EXU/CSRControl/_3291_ ( .A(\EXU/CSRControl/_0123_ ), .Z(\EXU/CSRControl/_1625_ ) );
BUF_X1 \EXU/CSRControl/_3292_ ( .A(\EXU/CSRControl/_0124_ ), .Z(\EXU/CSRControl/_1626_ ) );
BUF_X1 \EXU/CSRControl/_3293_ ( .A(\EXU/CSRControl/_0125_ ), .Z(\EXU/CSRControl/_1627_ ) );
BUF_X1 \EXU/CSRControl/_3294_ ( .A(\EXU/CSRControl/_0126_ ), .Z(\EXU/CSRControl/_1628_ ) );
BUF_X1 \EXU/CSRControl/_3295_ ( .A(\EXU/CSRControl/_0127_ ), .Z(\EXU/CSRControl/_1629_ ) );
BUF_X1 \EXU/CSRControl/_3296_ ( .A(\EXU/CSRControl/_0128_ ), .Z(\EXU/CSRControl/_1630_ ) );
BUF_X1 \EXU/CSRControl/_3297_ ( .A(\EXU/CSRControl/_0129_ ), .Z(\EXU/CSRControl/_1631_ ) );
BUF_X1 \EXU/CSRControl/_3298_ ( .A(\EXU/CSRControl/_0130_ ), .Z(\EXU/CSRControl/_1632_ ) );
BUF_X1 \EXU/CSRControl/_3299_ ( .A(\EXU/CSRControl/_0131_ ), .Z(\EXU/CSRControl/_1633_ ) );
INV_X1 \IDU/_011_ ( .A(\IDU/_000_ ), .ZN(\IDU/_009_ ) );
AND2_X1 \IDU/_012_ ( .A1(\IDU/_009_ ), .A2(\IDU/_005_ ), .ZN(\IDU/_001_ ) );
OR2_X4 \IDU/_013_ ( .A1(\IDU/_000_ ), .A2(\IDU/_006_ ), .ZN(\IDU/_002_ ) );
AND2_X1 \IDU/_014_ ( .A1(\IDU/_009_ ), .A2(\IDU/_007_ ), .ZN(\IDU/_003_ ) );
OR2_X4 \IDU/_015_ ( .A1(\IDU/_000_ ), .A2(\IDU/_008_ ), .ZN(\IDU/_004_ ) );
LOGIC0_X1 \IDU/_016_ ( .Z(\IDU/_010_ ) );
BUF_X1 \IDU/_017_ ( .A(\_IFU_io_out_bits_instruction [20] ), .Z(\_IDU_io_RegFileAccess_ra2 [0] ) );
BUF_X1 \IDU/_018_ ( .A(\_IFU_io_out_bits_instruction [21] ), .Z(\_IDU_io_RegFileAccess_ra2 [1] ) );
BUF_X1 \IDU/_019_ ( .A(\_IFU_io_out_bits_instruction [22] ), .Z(\_IDU_io_RegFileAccess_ra2 [2] ) );
BUF_X1 \IDU/_020_ ( .A(\_IFU_io_out_bits_instruction [23] ), .Z(\_IDU_io_RegFileAccess_ra2 [3] ) );
BUF_X1 \IDU/_021_ ( .A(_EXU_io_in_ready ), .Z(_IDU_io_in_ready ) );
BUF_X1 \IDU/_022_ ( .A(\_IFU_io_out_bits_pc [0] ), .Z(\_IDU_io_out_bits_pc [0] ) );
BUF_X1 \IDU/_023_ ( .A(\_IFU_io_out_bits_pc [1] ), .Z(\_IDU_io_out_bits_pc [1] ) );
BUF_X1 \IDU/_024_ ( .A(\_IFU_io_out_bits_pc [2] ), .Z(\_IDU_io_out_bits_pc [2] ) );
BUF_X1 \IDU/_025_ ( .A(\_IFU_io_out_bits_pc [3] ), .Z(\_IDU_io_out_bits_pc [3] ) );
BUF_X1 \IDU/_026_ ( .A(\_IFU_io_out_bits_pc [4] ), .Z(\_IDU_io_out_bits_pc [4] ) );
BUF_X1 \IDU/_027_ ( .A(\_IFU_io_out_bits_pc [5] ), .Z(\_IDU_io_out_bits_pc [5] ) );
BUF_X1 \IDU/_028_ ( .A(\_IFU_io_out_bits_pc [6] ), .Z(\_IDU_io_out_bits_pc [6] ) );
BUF_X1 \IDU/_029_ ( .A(\_IFU_io_out_bits_pc [7] ), .Z(\_IDU_io_out_bits_pc [7] ) );
BUF_X1 \IDU/_030_ ( .A(\_IFU_io_out_bits_pc [8] ), .Z(\_IDU_io_out_bits_pc [8] ) );
BUF_X1 \IDU/_031_ ( .A(\_IFU_io_out_bits_pc [9] ), .Z(\_IDU_io_out_bits_pc [9] ) );
BUF_X1 \IDU/_032_ ( .A(\_IFU_io_out_bits_pc [10] ), .Z(\_IDU_io_out_bits_pc [10] ) );
BUF_X1 \IDU/_033_ ( .A(\_IFU_io_out_bits_pc [11] ), .Z(\_IDU_io_out_bits_pc [11] ) );
BUF_X1 \IDU/_034_ ( .A(\_IFU_io_out_bits_pc [12] ), .Z(\_IDU_io_out_bits_pc [12] ) );
BUF_X1 \IDU/_035_ ( .A(\_IFU_io_out_bits_pc [13] ), .Z(\_IDU_io_out_bits_pc [13] ) );
BUF_X1 \IDU/_036_ ( .A(\_IFU_io_out_bits_pc [14] ), .Z(\_IDU_io_out_bits_pc [14] ) );
BUF_X1 \IDU/_037_ ( .A(\_IFU_io_out_bits_pc [15] ), .Z(\_IDU_io_out_bits_pc [15] ) );
BUF_X1 \IDU/_038_ ( .A(\_IFU_io_out_bits_pc [16] ), .Z(\_IDU_io_out_bits_pc [16] ) );
BUF_X1 \IDU/_039_ ( .A(\_IFU_io_out_bits_pc [17] ), .Z(\_IDU_io_out_bits_pc [17] ) );
BUF_X1 \IDU/_040_ ( .A(\_IFU_io_out_bits_pc [18] ), .Z(\_IDU_io_out_bits_pc [18] ) );
BUF_X1 \IDU/_041_ ( .A(\_IFU_io_out_bits_pc [19] ), .Z(\_IDU_io_out_bits_pc [19] ) );
BUF_X1 \IDU/_042_ ( .A(\_IFU_io_out_bits_pc [20] ), .Z(\_IDU_io_out_bits_pc [20] ) );
BUF_X1 \IDU/_043_ ( .A(\_IFU_io_out_bits_pc [21] ), .Z(\_IDU_io_out_bits_pc [21] ) );
BUF_X1 \IDU/_044_ ( .A(\_IFU_io_out_bits_pc [22] ), .Z(\_IDU_io_out_bits_pc [22] ) );
BUF_X1 \IDU/_045_ ( .A(\_IFU_io_out_bits_pc [23] ), .Z(\_IDU_io_out_bits_pc [23] ) );
BUF_X1 \IDU/_046_ ( .A(\_IFU_io_out_bits_pc [24] ), .Z(\_IDU_io_out_bits_pc [24] ) );
BUF_X1 \IDU/_047_ ( .A(\_IFU_io_out_bits_pc [25] ), .Z(\_IDU_io_out_bits_pc [25] ) );
BUF_X1 \IDU/_048_ ( .A(\_IFU_io_out_bits_pc [26] ), .Z(\_IDU_io_out_bits_pc [26] ) );
BUF_X1 \IDU/_049_ ( .A(\_IFU_io_out_bits_pc [27] ), .Z(\_IDU_io_out_bits_pc [27] ) );
BUF_X1 \IDU/_050_ ( .A(\_IFU_io_out_bits_pc [28] ), .Z(\_IDU_io_out_bits_pc [28] ) );
BUF_X1 \IDU/_051_ ( .A(\_IFU_io_out_bits_pc [29] ), .Z(\_IDU_io_out_bits_pc [29] ) );
BUF_X1 \IDU/_052_ ( .A(\_IFU_io_out_bits_pc [30] ), .Z(\_IDU_io_out_bits_pc [30] ) );
BUF_X1 \IDU/_053_ ( .A(\_IFU_io_out_bits_pc [31] ), .Z(\_IDU_io_out_bits_pc [31] ) );
BUF_X1 \IDU/_054_ ( .A(\_RegFile_io_rd1 [0] ), .Z(\_IDU_io_out_bits_rd1 [0] ) );
BUF_X1 \IDU/_055_ ( .A(\_RegFile_io_rd1 [1] ), .Z(\_IDU_io_out_bits_rd1 [1] ) );
BUF_X1 \IDU/_056_ ( .A(\_RegFile_io_rd1 [2] ), .Z(\_IDU_io_out_bits_rd1 [2] ) );
BUF_X1 \IDU/_057_ ( .A(\_RegFile_io_rd1 [3] ), .Z(\_IDU_io_out_bits_rd1 [3] ) );
BUF_X1 \IDU/_058_ ( .A(\_RegFile_io_rd1 [4] ), .Z(\_IDU_io_out_bits_rd1 [4] ) );
BUF_X1 \IDU/_059_ ( .A(\_RegFile_io_rd1 [5] ), .Z(\_IDU_io_out_bits_rd1 [5] ) );
BUF_X1 \IDU/_060_ ( .A(\_RegFile_io_rd1 [6] ), .Z(\_IDU_io_out_bits_rd1 [6] ) );
BUF_X1 \IDU/_061_ ( .A(\_RegFile_io_rd1 [7] ), .Z(\_IDU_io_out_bits_rd1 [7] ) );
BUF_X1 \IDU/_062_ ( .A(\_RegFile_io_rd1 [8] ), .Z(\_IDU_io_out_bits_rd1 [8] ) );
BUF_X1 \IDU/_063_ ( .A(\_RegFile_io_rd1 [9] ), .Z(\_IDU_io_out_bits_rd1 [9] ) );
BUF_X1 \IDU/_064_ ( .A(\_RegFile_io_rd1 [10] ), .Z(\_IDU_io_out_bits_rd1 [10] ) );
BUF_X1 \IDU/_065_ ( .A(\_RegFile_io_rd1 [11] ), .Z(\_IDU_io_out_bits_rd1 [11] ) );
BUF_X1 \IDU/_066_ ( .A(\_RegFile_io_rd1 [12] ), .Z(\_IDU_io_out_bits_rd1 [12] ) );
BUF_X1 \IDU/_067_ ( .A(\_RegFile_io_rd1 [13] ), .Z(\_IDU_io_out_bits_rd1 [13] ) );
BUF_X1 \IDU/_068_ ( .A(\_RegFile_io_rd1 [14] ), .Z(\_IDU_io_out_bits_rd1 [14] ) );
BUF_X1 \IDU/_069_ ( .A(\_RegFile_io_rd1 [15] ), .Z(\_IDU_io_out_bits_rd1 [15] ) );
BUF_X1 \IDU/_070_ ( .A(\_RegFile_io_rd1 [16] ), .Z(\_IDU_io_out_bits_rd1 [16] ) );
BUF_X1 \IDU/_071_ ( .A(\_RegFile_io_rd1 [17] ), .Z(\_IDU_io_out_bits_rd1 [17] ) );
BUF_X1 \IDU/_072_ ( .A(\_RegFile_io_rd1 [18] ), .Z(\_IDU_io_out_bits_rd1 [18] ) );
BUF_X1 \IDU/_073_ ( .A(\_RegFile_io_rd1 [19] ), .Z(\_IDU_io_out_bits_rd1 [19] ) );
BUF_X1 \IDU/_074_ ( .A(\_RegFile_io_rd1 [20] ), .Z(\_IDU_io_out_bits_rd1 [20] ) );
BUF_X1 \IDU/_075_ ( .A(\_RegFile_io_rd1 [21] ), .Z(\_IDU_io_out_bits_rd1 [21] ) );
BUF_X1 \IDU/_076_ ( .A(\_RegFile_io_rd1 [22] ), .Z(\_IDU_io_out_bits_rd1 [22] ) );
BUF_X1 \IDU/_077_ ( .A(\_RegFile_io_rd1 [23] ), .Z(\_IDU_io_out_bits_rd1 [23] ) );
BUF_X1 \IDU/_078_ ( .A(\_RegFile_io_rd1 [24] ), .Z(\_IDU_io_out_bits_rd1 [24] ) );
BUF_X1 \IDU/_079_ ( .A(\_RegFile_io_rd1 [25] ), .Z(\_IDU_io_out_bits_rd1 [25] ) );
BUF_X1 \IDU/_080_ ( .A(\_RegFile_io_rd1 [26] ), .Z(\_IDU_io_out_bits_rd1 [26] ) );
BUF_X1 \IDU/_081_ ( .A(\_RegFile_io_rd1 [27] ), .Z(\_IDU_io_out_bits_rd1 [27] ) );
BUF_X1 \IDU/_082_ ( .A(\_RegFile_io_rd1 [28] ), .Z(\_IDU_io_out_bits_rd1 [28] ) );
BUF_X1 \IDU/_083_ ( .A(\_RegFile_io_rd1 [29] ), .Z(\_IDU_io_out_bits_rd1 [29] ) );
BUF_X1 \IDU/_084_ ( .A(\_RegFile_io_rd1 [30] ), .Z(\_IDU_io_out_bits_rd1 [30] ) );
BUF_X1 \IDU/_085_ ( .A(\_RegFile_io_rd1 [31] ), .Z(\_IDU_io_out_bits_rd1 [31] ) );
BUF_X1 \IDU/_086_ ( .A(\_RegFile_io_rd2 [0] ), .Z(\_IDU_io_out_bits_rd2 [0] ) );
BUF_X1 \IDU/_087_ ( .A(\_RegFile_io_rd2 [1] ), .Z(\_IDU_io_out_bits_rd2 [1] ) );
BUF_X1 \IDU/_088_ ( .A(\_RegFile_io_rd2 [2] ), .Z(\_IDU_io_out_bits_rd2 [2] ) );
BUF_X1 \IDU/_089_ ( .A(\_RegFile_io_rd2 [3] ), .Z(\_IDU_io_out_bits_rd2 [3] ) );
BUF_X1 \IDU/_090_ ( .A(\_RegFile_io_rd2 [4] ), .Z(\_IDU_io_out_bits_rd2 [4] ) );
BUF_X1 \IDU/_091_ ( .A(\_RegFile_io_rd2 [5] ), .Z(\_IDU_io_out_bits_rd2 [5] ) );
BUF_X1 \IDU/_092_ ( .A(\_RegFile_io_rd2 [6] ), .Z(\_IDU_io_out_bits_rd2 [6] ) );
BUF_X1 \IDU/_093_ ( .A(\_RegFile_io_rd2 [7] ), .Z(\_IDU_io_out_bits_rd2 [7] ) );
BUF_X1 \IDU/_094_ ( .A(\_RegFile_io_rd2 [8] ), .Z(\_IDU_io_out_bits_rd2 [8] ) );
BUF_X1 \IDU/_095_ ( .A(\_RegFile_io_rd2 [9] ), .Z(\_IDU_io_out_bits_rd2 [9] ) );
BUF_X1 \IDU/_096_ ( .A(\_RegFile_io_rd2 [10] ), .Z(\_IDU_io_out_bits_rd2 [10] ) );
BUF_X1 \IDU/_097_ ( .A(\_RegFile_io_rd2 [11] ), .Z(\_IDU_io_out_bits_rd2 [11] ) );
BUF_X1 \IDU/_098_ ( .A(\_RegFile_io_rd2 [12] ), .Z(\_IDU_io_out_bits_rd2 [12] ) );
BUF_X1 \IDU/_099_ ( .A(\_RegFile_io_rd2 [13] ), .Z(\_IDU_io_out_bits_rd2 [13] ) );
BUF_X1 \IDU/_100_ ( .A(\_RegFile_io_rd2 [14] ), .Z(\_IDU_io_out_bits_rd2 [14] ) );
BUF_X1 \IDU/_101_ ( .A(\_RegFile_io_rd2 [15] ), .Z(\_IDU_io_out_bits_rd2 [15] ) );
BUF_X1 \IDU/_102_ ( .A(\_RegFile_io_rd2 [16] ), .Z(\_IDU_io_out_bits_rd2 [16] ) );
BUF_X1 \IDU/_103_ ( .A(\_RegFile_io_rd2 [17] ), .Z(\_IDU_io_out_bits_rd2 [17] ) );
BUF_X1 \IDU/_104_ ( .A(\_RegFile_io_rd2 [18] ), .Z(\_IDU_io_out_bits_rd2 [18] ) );
BUF_X1 \IDU/_105_ ( .A(\_RegFile_io_rd2 [19] ), .Z(\_IDU_io_out_bits_rd2 [19] ) );
BUF_X1 \IDU/_106_ ( .A(\_RegFile_io_rd2 [20] ), .Z(\_IDU_io_out_bits_rd2 [20] ) );
BUF_X1 \IDU/_107_ ( .A(\_RegFile_io_rd2 [21] ), .Z(\_IDU_io_out_bits_rd2 [21] ) );
BUF_X1 \IDU/_108_ ( .A(\_RegFile_io_rd2 [22] ), .Z(\_IDU_io_out_bits_rd2 [22] ) );
BUF_X1 \IDU/_109_ ( .A(\_RegFile_io_rd2 [23] ), .Z(\_IDU_io_out_bits_rd2 [23] ) );
BUF_X1 \IDU/_110_ ( .A(\_RegFile_io_rd2 [24] ), .Z(\_IDU_io_out_bits_rd2 [24] ) );
BUF_X1 \IDU/_111_ ( .A(\_RegFile_io_rd2 [25] ), .Z(\_IDU_io_out_bits_rd2 [25] ) );
BUF_X1 \IDU/_112_ ( .A(\_RegFile_io_rd2 [26] ), .Z(\_IDU_io_out_bits_rd2 [26] ) );
BUF_X1 \IDU/_113_ ( .A(\_RegFile_io_rd2 [27] ), .Z(\_IDU_io_out_bits_rd2 [27] ) );
BUF_X1 \IDU/_114_ ( .A(\_RegFile_io_rd2 [28] ), .Z(\_IDU_io_out_bits_rd2 [28] ) );
BUF_X1 \IDU/_115_ ( .A(\_RegFile_io_rd2 [29] ), .Z(\_IDU_io_out_bits_rd2 [29] ) );
BUF_X1 \IDU/_116_ ( .A(\_RegFile_io_rd2 [30] ), .Z(\_IDU_io_out_bits_rd2 [30] ) );
BUF_X1 \IDU/_117_ ( .A(\_RegFile_io_rd2 [31] ), .Z(\_IDU_io_out_bits_rd2 [31] ) );
BUF_X1 \IDU/_118_ ( .A(\_IFU_io_out_bits_instruction [15] ), .Z(\_IDU_io_out_bits_uimm [0] ) );
BUF_X1 \IDU/_119_ ( .A(\_IFU_io_out_bits_instruction [16] ), .Z(\_IDU_io_out_bits_uimm [1] ) );
BUF_X1 \IDU/_120_ ( .A(\_IFU_io_out_bits_instruction [17] ), .Z(\_IDU_io_out_bits_uimm [2] ) );
BUF_X1 \IDU/_121_ ( .A(\_IFU_io_out_bits_instruction [18] ), .Z(\_IDU_io_out_bits_uimm [3] ) );
BUF_X1 \IDU/_122_ ( .A(\_IFU_io_out_bits_instruction [19] ), .Z(\_IDU_io_out_bits_uimm [4] ) );
BUF_X1 \IDU/_123_ ( .A(\IDU/_010_ ), .Z(\_IDU_io_out_bits_uimm [5] ) );
BUF_X1 \IDU/_124_ ( .A(\IDU/_010_ ), .Z(\_IDU_io_out_bits_uimm [6] ) );
BUF_X1 \IDU/_125_ ( .A(\IDU/_010_ ), .Z(\_IDU_io_out_bits_uimm [7] ) );
BUF_X1 \IDU/_126_ ( .A(\IDU/_010_ ), .Z(\_IDU_io_out_bits_uimm [8] ) );
BUF_X1 \IDU/_127_ ( .A(\IDU/_010_ ), .Z(\_IDU_io_out_bits_uimm [9] ) );
BUF_X1 \IDU/_128_ ( .A(\IDU/_010_ ), .Z(\_IDU_io_out_bits_uimm [10] ) );
BUF_X1 \IDU/_129_ ( .A(\IDU/_010_ ), .Z(\_IDU_io_out_bits_uimm [11] ) );
BUF_X1 \IDU/_130_ ( .A(\IDU/_010_ ), .Z(\_IDU_io_out_bits_uimm [12] ) );
BUF_X1 \IDU/_131_ ( .A(\IDU/_010_ ), .Z(\_IDU_io_out_bits_uimm [13] ) );
BUF_X1 \IDU/_132_ ( .A(\IDU/_010_ ), .Z(\_IDU_io_out_bits_uimm [14] ) );
BUF_X1 \IDU/_133_ ( .A(\IDU/_010_ ), .Z(\_IDU_io_out_bits_uimm [15] ) );
BUF_X1 \IDU/_134_ ( .A(\IDU/_010_ ), .Z(\_IDU_io_out_bits_uimm [16] ) );
BUF_X1 \IDU/_135_ ( .A(\IDU/_010_ ), .Z(\_IDU_io_out_bits_uimm [17] ) );
BUF_X1 \IDU/_136_ ( .A(\IDU/_010_ ), .Z(\_IDU_io_out_bits_uimm [18] ) );
BUF_X1 \IDU/_137_ ( .A(\IDU/_010_ ), .Z(\_IDU_io_out_bits_uimm [19] ) );
BUF_X1 \IDU/_138_ ( .A(\IDU/_010_ ), .Z(\_IDU_io_out_bits_uimm [20] ) );
BUF_X1 \IDU/_139_ ( .A(\IDU/_010_ ), .Z(\_IDU_io_out_bits_uimm [21] ) );
BUF_X1 \IDU/_140_ ( .A(\IDU/_010_ ), .Z(\_IDU_io_out_bits_uimm [22] ) );
BUF_X1 \IDU/_141_ ( .A(\IDU/_010_ ), .Z(\_IDU_io_out_bits_uimm [23] ) );
BUF_X1 \IDU/_142_ ( .A(\IDU/_010_ ), .Z(\_IDU_io_out_bits_uimm [24] ) );
BUF_X1 \IDU/_143_ ( .A(\IDU/_010_ ), .Z(\_IDU_io_out_bits_uimm [25] ) );
BUF_X1 \IDU/_144_ ( .A(\IDU/_010_ ), .Z(\_IDU_io_out_bits_uimm [26] ) );
BUF_X1 \IDU/_145_ ( .A(\IDU/_010_ ), .Z(\_IDU_io_out_bits_uimm [27] ) );
BUF_X1 \IDU/_146_ ( .A(\IDU/_010_ ), .Z(\_IDU_io_out_bits_uimm [28] ) );
BUF_X1 \IDU/_147_ ( .A(\IDU/_010_ ), .Z(\_IDU_io_out_bits_uimm [29] ) );
BUF_X1 \IDU/_148_ ( .A(\IDU/_010_ ), .Z(\_IDU_io_out_bits_uimm [30] ) );
BUF_X1 \IDU/_149_ ( .A(\IDU/_010_ ), .Z(\_IDU_io_out_bits_uimm [31] ) );
BUF_X1 \IDU/_150_ ( .A(\_IFU_io_out_bits_instruction [7] ), .Z(\_IDU_io_out_bits_wa [0] ) );
BUF_X1 \IDU/_151_ ( .A(\_IFU_io_out_bits_instruction [8] ), .Z(\_IDU_io_out_bits_wa [1] ) );
BUF_X1 \IDU/_152_ ( .A(\_IFU_io_out_bits_instruction [9] ), .Z(\_IDU_io_out_bits_wa [2] ) );
BUF_X1 \IDU/_153_ ( .A(\_IFU_io_out_bits_instruction [10] ), .Z(\_IDU_io_out_bits_wa [3] ) );
BUF_X1 \IDU/_154_ ( .A(\_IFU_io_out_bits_instruction [11] ), .Z(\_IDU_io_out_bits_wa [4] ) );
BUF_X1 \IDU/_155_ ( .A(_IFU_io_out_valid ), .Z(_IDU_io_out_valid ) );
BUF_X1 \IDU/_156_ ( .A(\_IFU_io_out_bits_instruction [15] ), .Z(\IDU/_005_ ) );
BUF_X1 \IDU/_157_ ( .A(\IDU/_Control_io_isEnd ), .Z(\IDU/_000_ ) );
BUF_X1 \IDU/_158_ ( .A(\IDU/_001_ ), .Z(\_IDU_io_RegFileAccess_ra1 [0] ) );
BUF_X1 \IDU/_159_ ( .A(\_IFU_io_out_bits_instruction [16] ), .Z(\IDU/_006_ ) );
BUF_X1 \IDU/_160_ ( .A(\IDU/_002_ ), .Z(\_IDU_io_RegFileAccess_ra1 [1] ) );
BUF_X1 \IDU/_161_ ( .A(\_IFU_io_out_bits_instruction [17] ), .Z(\IDU/_007_ ) );
BUF_X1 \IDU/_162_ ( .A(\IDU/_003_ ), .Z(\_IDU_io_RegFileAccess_ra1 [2] ) );
BUF_X1 \IDU/_163_ ( .A(\_IFU_io_out_bits_instruction [18] ), .Z(\IDU/_008_ ) );
BUF_X1 \IDU/_164_ ( .A(\IDU/_004_ ), .Z(\_IDU_io_RegFileAccess_ra1 [3] ) );
AND2_X1 \IDU/Control/_121_ ( .A1(\IDU/Control/_042_ ), .A2(\IDU/Control/_038_ ), .ZN(\IDU/Control/_082_ ) );
NAND2_X1 \IDU/Control/_122_ ( .A1(\IDU/Control/_082_ ), .A2(\IDU/Control/_043_ ), .ZN(\IDU/Control/_083_ ) );
INV_X4 \IDU/Control/_123_ ( .A(\IDU/Control/_038_ ), .ZN(\IDU/Control/_084_ ) );
INV_X32 \IDU/Control/_124_ ( .A(\IDU/Control/_020_ ), .ZN(\IDU/Control/_085_ ) );
NAND4_X1 \IDU/Control/_125_ ( .A1(\IDU/Control/_084_ ), .A2(\IDU/Control/_085_ ), .A3(\IDU/Control/_019_ ), .A4(\IDU/Control/_042_ ), .ZN(\IDU/Control/_086_ ) );
NAND4_X1 \IDU/Control/_126_ ( .A1(\IDU/Control/_084_ ), .A2(\IDU/Control/_019_ ), .A3(\IDU/Control/_042_ ), .A4(\IDU/Control/_021_ ), .ZN(\IDU/Control/_087_ ) );
NAND3_X1 \IDU/Control/_127_ ( .A1(\IDU/Control/_083_ ), .A2(\IDU/Control/_086_ ), .A3(\IDU/Control/_087_ ), .ZN(\IDU/Control/_003_ ) );
AND2_X1 \IDU/Control/_128_ ( .A1(\IDU/Control/_084_ ), .A2(\IDU/Control/_021_ ), .ZN(\IDU/Control/_088_ ) );
INV_X1 \IDU/Control/_129_ ( .A(\IDU/Control/_043_ ), .ZN(\IDU/Control/_089_ ) );
NOR2_X1 \IDU/Control/_130_ ( .A1(\IDU/Control/_089_ ), .A2(\IDU/Control/_042_ ), .ZN(\IDU/Control/_090_ ) );
NAND2_X1 \IDU/Control/_131_ ( .A1(\IDU/Control/_088_ ), .A2(\IDU/Control/_090_ ), .ZN(\IDU/Control/_091_ ) );
NAND3_X1 \IDU/Control/_132_ ( .A1(\IDU/Control/_084_ ), .A2(\IDU/Control/_042_ ), .A3(\IDU/Control/_020_ ), .ZN(\IDU/Control/_092_ ) );
NAND3_X1 \IDU/Control/_133_ ( .A1(\IDU/Control/_091_ ), .A2(\IDU/Control/_083_ ), .A3(\IDU/Control/_092_ ), .ZN(\IDU/Control/_004_ ) );
AND3_X1 \IDU/Control/_134_ ( .A1(\IDU/Control/_084_ ), .A2(\IDU/Control/_042_ ), .A3(\IDU/Control/_021_ ), .ZN(\IDU/Control/_012_ ) );
AND3_X1 \IDU/Control/_135_ ( .A1(\IDU/Control/_084_ ), .A2(\IDU/Control/_019_ ), .A3(\IDU/Control/_042_ ), .ZN(\IDU/Control/_093_ ) );
AND2_X1 \IDU/Control/_136_ ( .A1(\IDU/Control/_042_ ), .A2(\IDU/Control/_043_ ), .ZN(\IDU/Control/_094_ ) );
OAI21_X1 \IDU/Control/_137_ ( .A(\IDU/Control/_039_ ), .B1(\IDU/Control/_093_ ), .B2(\IDU/Control/_094_ ), .ZN(\IDU/Control/_095_ ) );
INV_X32 \IDU/Control/_138_ ( .A(\IDU/Control/_044_ ), .ZN(\IDU/Control/_096_ ) );
NOR3_X1 \IDU/Control/_139_ ( .A1(\IDU/Control/_096_ ), .A2(\IDU/Control/_038_ ), .A3(\IDU/Control/_021_ ), .ZN(\IDU/Control/_097_ ) );
INV_X16 \IDU/Control/_140_ ( .A(\IDU/Control/_042_ ), .ZN(\IDU/Control/_098_ ) );
NAND2_X1 \IDU/Control/_141_ ( .A1(\IDU/Control/_097_ ), .A2(\IDU/Control/_098_ ), .ZN(\IDU/Control/_099_ ) );
NOR2_X1 \IDU/Control/_142_ ( .A1(\IDU/Control/_085_ ), .A2(\IDU/Control/_038_ ), .ZN(\IDU/Control/_100_ ) );
OAI21_X1 \IDU/Control/_143_ ( .A(\IDU/Control/_100_ ), .B1(\IDU/Control/_019_ ), .B2(\IDU/Control/_044_ ), .ZN(\IDU/Control/_101_ ) );
NAND3_X1 \IDU/Control/_144_ ( .A1(\IDU/Control/_095_ ), .A2(\IDU/Control/_099_ ), .A3(\IDU/Control/_101_ ), .ZN(\IDU/Control/_005_ ) );
INV_X4 \IDU/Control/_145_ ( .A(\IDU/Control/_019_ ), .ZN(\IDU/Control/_102_ ) );
NOR2_X1 \IDU/Control/_146_ ( .A1(\IDU/Control/_102_ ), .A2(\IDU/Control/_038_ ), .ZN(\IDU/Control/_103_ ) );
AND2_X4 \IDU/Control/_147_ ( .A1(\IDU/Control/_027_ ), .A2(\IDU/Control/_016_ ), .ZN(\IDU/Control/_104_ ) );
AND3_X1 \IDU/Control/_148_ ( .A1(\IDU/Control/_103_ ), .A2(\IDU/Control/_094_ ), .A3(\IDU/Control/_104_ ), .ZN(\IDU/Control/_105_ ) );
NOR2_X1 \IDU/Control/_149_ ( .A1(\IDU/Control/_096_ ), .A2(\IDU/Control/_041_ ), .ZN(\IDU/Control/_106_ ) );
NAND2_X1 \IDU/Control/_150_ ( .A1(\IDU/Control/_105_ ), .A2(\IDU/Control/_106_ ), .ZN(\IDU/Control/_107_ ) );
NOR4_X4 \IDU/Control/_151_ ( .A1(\IDU/Control/_028_ ), .A2(\IDU/Control/_031_ ), .A3(\IDU/Control/_030_ ), .A4(\IDU/Control/_033_ ), .ZN(\IDU/Control/_108_ ) );
NOR4_X4 \IDU/Control/_152_ ( .A1(\IDU/Control/_039_ ), .A2(\IDU/Control/_023_ ), .A3(\IDU/Control/_022_ ), .A4(\IDU/Control/_024_ ), .ZN(\IDU/Control/_109_ ) );
AND2_X2 \IDU/Control/_153_ ( .A1(\IDU/Control/_108_ ), .A2(\IDU/Control/_109_ ), .ZN(\IDU/Control/_110_ ) );
AND2_X1 \IDU/Control/_154_ ( .A1(\IDU/Control/_094_ ), .A2(\IDU/Control/_104_ ), .ZN(\IDU/Control/_111_ ) );
NOR4_X4 \IDU/Control/_155_ ( .A1(\IDU/Control/_032_ ), .A2(\IDU/Control/_035_ ), .A3(\IDU/Control/_034_ ), .A4(\IDU/Control/_040_ ), .ZN(\IDU/Control/_112_ ) );
NAND3_X2 \IDU/Control/_156_ ( .A1(\IDU/Control/_110_ ), .A2(\IDU/Control/_111_ ), .A3(\IDU/Control/_112_ ), .ZN(\IDU/Control/_113_ ) );
AND4_X2 \IDU/Control/_157_ ( .A1(\IDU/Control/_102_ ), .A2(\IDU/Control/_084_ ), .A3(\IDU/Control/_085_ ), .A4(\IDU/Control/_044_ ), .ZN(\IDU/Control/_114_ ) );
INV_X1 \IDU/Control/_158_ ( .A(\IDU/Control/_046_ ), .ZN(\IDU/Control/_115_ ) );
AND4_X1 \IDU/Control/_159_ ( .A1(\IDU/Control/_029_ ), .A2(\IDU/Control/_115_ ), .A3(\IDU/Control/_037_ ), .A4(\IDU/Control/_036_ ), .ZN(\IDU/Control/_116_ ) );
AND2_X1 \IDU/Control/_160_ ( .A1(\IDU/Control/_114_ ), .A2(\IDU/Control/_116_ ), .ZN(\IDU/Control/_117_ ) );
NOR4_X1 \IDU/Control/_161_ ( .A1(\IDU/Control/_021_ ), .A2(\IDU/Control/_041_ ), .A3(\IDU/Control/_017_ ), .A4(\IDU/Control/_018_ ), .ZN(\IDU/Control/_118_ ) );
NOR4_X1 \IDU/Control/_162_ ( .A1(\IDU/Control/_045_ ), .A2(\IDU/Control/_047_ ), .A3(\IDU/Control/_025_ ), .A4(\IDU/Control/_026_ ), .ZN(\IDU/Control/_119_ ) );
NAND3_X1 \IDU/Control/_163_ ( .A1(\IDU/Control/_117_ ), .A2(\IDU/Control/_118_ ), .A3(\IDU/Control/_119_ ), .ZN(\IDU/Control/_120_ ) );
OAI21_X1 \IDU/Control/_164_ ( .A(\IDU/Control/_107_ ), .B1(\IDU/Control/_113_ ), .B2(\IDU/Control/_120_ ), .ZN(\IDU/Control/_009_ ) );
AND4_X1 \IDU/Control/_165_ ( .A1(\IDU/Control/_094_ ), .A2(\IDU/Control/_100_ ), .A3(\IDU/Control/_106_ ), .A4(\IDU/Control/_104_ ), .ZN(\IDU/Control/_010_ ) );
NOR4_X1 \IDU/Control/_166_ ( .A1(\IDU/Control/_021_ ), .A2(\IDU/Control/_041_ ), .A3(\IDU/Control/_045_ ), .A4(\IDU/Control/_047_ ), .ZN(\IDU/Control/_054_ ) );
NOR4_X1 \IDU/Control/_167_ ( .A1(\IDU/Control/_019_ ), .A2(\IDU/Control/_020_ ), .A3(\IDU/Control/_025_ ), .A4(\IDU/Control/_026_ ), .ZN(\IDU/Control/_055_ ) );
NOR4_X1 \IDU/Control/_168_ ( .A1(\IDU/Control/_029_ ), .A2(\IDU/Control/_037_ ), .A3(\IDU/Control/_036_ ), .A4(\IDU/Control/_046_ ), .ZN(\IDU/Control/_056_ ) );
NOR4_X1 \IDU/Control/_169_ ( .A1(\IDU/Control/_096_ ), .A2(\IDU/Control/_038_ ), .A3(\IDU/Control/_017_ ), .A4(\IDU/Control/_018_ ), .ZN(\IDU/Control/_057_ ) );
NAND4_X1 \IDU/Control/_170_ ( .A1(\IDU/Control/_054_ ), .A2(\IDU/Control/_055_ ), .A3(\IDU/Control/_056_ ), .A4(\IDU/Control/_057_ ), .ZN(\IDU/Control/_058_ ) );
AOI21_X1 \IDU/Control/_171_ ( .A(\IDU/Control/_113_ ), .B1(\IDU/Control/_120_ ), .B2(\IDU/Control/_058_ ), .ZN(\IDU/Control/_011_ ) );
AND2_X4 \IDU/Control/_172_ ( .A1(\IDU/Control/_043_ ), .A2(\IDU/Control/_044_ ), .ZN(\IDU/Control/_059_ ) );
AND2_X2 \IDU/Control/_173_ ( .A1(\IDU/Control/_104_ ), .A2(\IDU/Control/_059_ ), .ZN(\IDU/Control/_060_ ) );
INV_X1 \IDU/Control/_174_ ( .A(\IDU/Control/_041_ ), .ZN(\IDU/Control/_061_ ) );
AND3_X4 \IDU/Control/_175_ ( .A1(\IDU/Control/_060_ ), .A2(\IDU/Control/_098_ ), .A3(\IDU/Control/_061_ ), .ZN(\IDU/Control/_062_ ) );
NAND3_X2 \IDU/Control/_176_ ( .A1(\IDU/Control/_062_ ), .A2(\IDU/Control/_085_ ), .A3(\IDU/Control/_103_ ), .ZN(\IDU/Control/_063_ ) );
AND3_X1 \IDU/Control/_177_ ( .A1(\IDU/Control/_098_ ), .A2(\IDU/Control/_043_ ), .A3(\IDU/Control/_044_ ), .ZN(\IDU/Control/_064_ ) );
AND4_X1 \IDU/Control/_178_ ( .A1(\IDU/Control/_038_ ), .A2(\IDU/Control/_027_ ), .A3(\IDU/Control/_016_ ), .A4(\IDU/Control/_041_ ), .ZN(\IDU/Control/_065_ ) );
NAND2_X1 \IDU/Control/_179_ ( .A1(\IDU/Control/_064_ ), .A2(\IDU/Control/_065_ ), .ZN(\IDU/Control/_066_ ) );
NOR2_X1 \IDU/Control/_180_ ( .A1(\IDU/Control/_038_ ), .A2(\IDU/Control/_041_ ), .ZN(\IDU/Control/_067_ ) );
NAND4_X1 \IDU/Control/_181_ ( .A1(\IDU/Control/_060_ ), .A2(\IDU/Control/_019_ ), .A3(\IDU/Control/_021_ ), .A4(\IDU/Control/_067_ ), .ZN(\IDU/Control/_068_ ) );
OAI211_X2 \IDU/Control/_182_ ( .A(\IDU/Control/_063_ ), .B(\IDU/Control/_066_ ), .C1(\IDU/Control/_042_ ), .C2(\IDU/Control/_068_ ), .ZN(\IDU/Control/_006_ ) );
NAND2_X1 \IDU/Control/_183_ ( .A1(\IDU/Control/_062_ ), .A2(\IDU/Control/_088_ ), .ZN(\IDU/Control/_069_ ) );
NOR4_X1 \IDU/Control/_184_ ( .A1(\IDU/Control/_096_ ), .A2(\IDU/Control/_021_ ), .A3(\IDU/Control/_020_ ), .A4(\IDU/Control/_041_ ), .ZN(\IDU/Control/_070_ ) );
AND4_X1 \IDU/Control/_185_ ( .A1(\IDU/Control/_102_ ), .A2(\IDU/Control/_098_ ), .A3(\IDU/Control/_038_ ), .A4(\IDU/Control/_043_ ), .ZN(\IDU/Control/_071_ ) );
NAND3_X1 \IDU/Control/_186_ ( .A1(\IDU/Control/_070_ ), .A2(\IDU/Control/_071_ ), .A3(\IDU/Control/_104_ ), .ZN(\IDU/Control/_072_ ) );
NAND2_X1 \IDU/Control/_187_ ( .A1(\IDU/Control/_069_ ), .A2(\IDU/Control/_072_ ), .ZN(\IDU/Control/_007_ ) );
NAND4_X1 \IDU/Control/_188_ ( .A1(\IDU/Control/_060_ ), .A2(\IDU/Control/_098_ ), .A3(\IDU/Control/_085_ ), .A4(\IDU/Control/_067_ ), .ZN(\IDU/Control/_073_ ) );
NAND2_X1 \IDU/Control/_189_ ( .A1(\IDU/Control/_069_ ), .A2(\IDU/Control/_073_ ), .ZN(\IDU/Control/_008_ ) );
NAND2_X1 \IDU/Control/_190_ ( .A1(\IDU/Control/_042_ ), .A2(\IDU/Control/_044_ ), .ZN(\IDU/Control/_074_ ) );
NOR4_X1 \IDU/Control/_191_ ( .A1(\IDU/Control/_074_ ), .A2(\IDU/Control/_019_ ), .A3(\IDU/Control/_020_ ), .A4(\IDU/Control/_028_ ), .ZN(\IDU/Control/_051_ ) );
AND3_X1 \IDU/Control/_192_ ( .A1(\IDU/Control/_104_ ), .A2(\IDU/Control/_089_ ), .A3(\IDU/Control/_096_ ), .ZN(\IDU/Control/_075_ ) );
OAI21_X1 \IDU/Control/_193_ ( .A(\IDU/Control/_020_ ), .B1(\IDU/Control/_019_ ), .B2(\IDU/Control/_021_ ), .ZN(\IDU/Control/_076_ ) );
AND4_X1 \IDU/Control/_194_ ( .A1(\IDU/Control/_098_ ), .A2(\IDU/Control/_075_ ), .A3(\IDU/Control/_067_ ), .A4(\IDU/Control/_076_ ), .ZN(\IDU/Control/_049_ ) );
INV_X1 \IDU/Control/_195_ ( .A(\IDU/Control/_010_ ), .ZN(\IDU/Control/_077_ ) );
NAND2_X1 \IDU/Control/_196_ ( .A1(\IDU/Control/_077_ ), .A2(\IDU/Control/_107_ ), .ZN(\IDU/Control/_053_ ) );
NAND4_X1 \IDU/Control/_197_ ( .A1(\IDU/Control/_102_ ), .A2(\IDU/Control/_042_ ), .A3(\IDU/Control/_044_ ), .A4(\IDU/Control/_028_ ), .ZN(\IDU/Control/_078_ ) );
NOR2_X1 \IDU/Control/_198_ ( .A1(\IDU/Control/_078_ ), .A2(\IDU/Control/_020_ ), .ZN(\IDU/Control/_048_ ) );
INV_X1 \IDU/Control/_199_ ( .A(\IDU/Control/_082_ ), .ZN(\IDU/Control/_079_ ) );
NAND3_X1 \IDU/Control/_200_ ( .A1(\IDU/Control/_099_ ), .A2(\IDU/Control/_091_ ), .A3(\IDU/Control/_079_ ), .ZN(\IDU/Control/_013_ ) );
AND2_X1 \IDU/Control/_201_ ( .A1(\IDU/Control/_090_ ), .A2(\IDU/Control/_096_ ), .ZN(\IDU/Control/_050_ ) );
INV_X1 \IDU/Control/_202_ ( .A(\IDU/Control/_050_ ), .ZN(\IDU/Control/_080_ ) );
NAND3_X1 \IDU/Control/_203_ ( .A1(\IDU/Control/_080_ ), .A2(\IDU/Control/_091_ ), .A3(\IDU/Control/_099_ ), .ZN(\IDU/Control/_014_ ) );
AND2_X1 \IDU/Control/_204_ ( .A1(\IDU/Control/_043_ ), .A2(\IDU/Control/_041_ ), .ZN(\IDU/Control/_015_ ) );
AND2_X1 \IDU/Control/_205_ ( .A1(\IDU/Control/_038_ ), .A2(\IDU/Control/_044_ ), .ZN(\IDU/Control/_002_ ) );
OAI211_X2 \IDU/Control/_206_ ( .A(\IDU/Control/_098_ ), .B(\IDU/Control/_043_ ), .C1(\IDU/Control/_084_ ), .C2(\IDU/Control/_096_ ), .ZN(\IDU/Control/_052_ ) );
NAND3_X1 \IDU/Control/_207_ ( .A1(\IDU/Control/_075_ ), .A2(\IDU/Control/_061_ ), .A3(\IDU/Control/_082_ ), .ZN(\IDU/Control/_081_ ) );
NAND3_X1 \IDU/Control/_208_ ( .A1(\IDU/Control/_081_ ), .A2(\IDU/Control/_066_ ), .A3(\IDU/Control/_072_ ), .ZN(\IDU/Control/_000_ ) );
NAND4_X1 \IDU/Control/_209_ ( .A1(\IDU/Control/_080_ ), .A2(\IDU/Control/_043_ ), .A3(\IDU/Control/_079_ ), .A4(\IDU/Control/_074_ ), .ZN(\IDU/Control/_001_ ) );
BUF_X1 \IDU/Control/_210_ ( .A(_IDU_io_out_bits_control_csrSrc ), .Z(\_IDU_io_out_bits_control_aluCtr [2] ) );
BUF_X1 \IDU/Control/_211_ ( .A(\_IFU_io_out_bits_instruction [12] ), .Z(\_IDU_io_out_bits_control_memOp [0] ) );
BUF_X1 \IDU/Control/_212_ ( .A(\_IFU_io_out_bits_instruction [13] ), .Z(\_IDU_io_out_bits_control_memOp [1] ) );
BUF_X1 \IDU/Control/_213_ ( .A(\_IFU_io_out_bits_instruction [14] ), .Z(\_IDU_io_out_bits_control_memOp [2] ) );
BUF_X1 \IDU/Control/_214_ ( .A(_IDU_io_out_bits_control_memRen ), .Z(\_IDU_io_out_bits_control_wbSrc [0] ) );
BUF_X1 \IDU/Control/_215_ ( .A(\_IFU_io_out_bits_instruction [12] ), .Z(\IDU/Control/_019_ ) );
BUF_X1 \IDU/Control/_216_ ( .A(\_IFU_io_out_bits_instruction [4] ), .Z(\IDU/Control/_042_ ) );
BUF_X1 \IDU/Control/_217_ ( .A(\_IFU_io_out_bits_instruction [2] ), .Z(\IDU/Control/_038_ ) );
BUF_X1 \IDU/Control/_218_ ( .A(\_IFU_io_out_bits_instruction [14] ), .Z(\IDU/Control/_021_ ) );
BUF_X1 \IDU/Control/_219_ ( .A(\_IFU_io_out_bits_instruction [13] ), .Z(\IDU/Control/_020_ ) );
BUF_X1 \IDU/Control/_220_ ( .A(\_IFU_io_out_bits_instruction [5] ), .Z(\IDU/Control/_043_ ) );
BUF_X1 \IDU/Control/_221_ ( .A(\IDU/Control/_003_ ), .Z(\_IDU_io_out_bits_control_aluCtr [0] ) );
BUF_X1 \IDU/Control/_222_ ( .A(\IDU/Control/_004_ ), .Z(\_IDU_io_out_bits_control_aluCtr [1] ) );
BUF_X1 \IDU/Control/_223_ ( .A(\IDU/Control/_012_ ), .Z(_IDU_io_out_bits_control_csrSrc ) );
BUF_X1 \IDU/Control/_224_ ( .A(\_IFU_io_out_bits_instruction [6] ), .Z(\IDU/Control/_044_ ) );
BUF_X1 \IDU/Control/_225_ ( .A(\_IFU_io_out_bits_instruction [30] ), .Z(\IDU/Control/_039_ ) );
BUF_X1 \IDU/Control/_226_ ( .A(\IDU/Control/_005_ ), .Z(\_IDU_io_out_bits_control_aluCtr [3] ) );
BUF_X1 \IDU/Control/_227_ ( .A(\_IFU_io_out_bits_instruction [1] ), .Z(\IDU/Control/_027_ ) );
BUF_X1 \IDU/Control/_228_ ( .A(\_IFU_io_out_bits_instruction [0] ), .Z(\IDU/Control/_016_ ) );
BUF_X1 \IDU/Control/_229_ ( .A(\_IFU_io_out_bits_instruction [3] ), .Z(\IDU/Control/_041_ ) );
BUF_X1 \IDU/Control/_230_ ( .A(\_IFU_io_out_bits_instruction [21] ), .Z(\IDU/Control/_029_ ) );
BUF_X1 \IDU/Control/_231_ ( .A(\_IFU_io_out_bits_instruction [29] ), .Z(\IDU/Control/_037_ ) );
BUF_X1 \IDU/Control/_232_ ( .A(\_IFU_io_out_bits_instruction [28] ), .Z(\IDU/Control/_036_ ) );
BUF_X1 \IDU/Control/_233_ ( .A(\_IFU_io_out_bits_instruction [8] ), .Z(\IDU/Control/_046_ ) );
BUF_X1 \IDU/Control/_234_ ( .A(\_IFU_io_out_bits_instruction [7] ), .Z(\IDU/Control/_045_ ) );
BUF_X1 \IDU/Control/_235_ ( .A(\_IFU_io_out_bits_instruction [10] ), .Z(\IDU/Control/_017_ ) );
BUF_X1 \IDU/Control/_236_ ( .A(\_IFU_io_out_bits_instruction [9] ), .Z(\IDU/Control/_047_ ) );
BUF_X1 \IDU/Control/_237_ ( .A(\_IFU_io_out_bits_instruction [11] ), .Z(\IDU/Control/_018_ ) );
BUF_X1 \IDU/Control/_238_ ( .A(\_IFU_io_out_bits_instruction [16] ), .Z(\IDU/Control/_023_ ) );
BUF_X1 \IDU/Control/_239_ ( .A(\_IFU_io_out_bits_instruction [15] ), .Z(\IDU/Control/_022_ ) );
BUF_X1 \IDU/Control/_240_ ( .A(\_IFU_io_out_bits_instruction [18] ), .Z(\IDU/Control/_025_ ) );
BUF_X1 \IDU/Control/_241_ ( .A(\_IFU_io_out_bits_instruction [17] ), .Z(\IDU/Control/_024_ ) );
BUF_X1 \IDU/Control/_242_ ( .A(\_IFU_io_out_bits_instruction [19] ), .Z(\IDU/Control/_026_ ) );
BUF_X1 \IDU/Control/_243_ ( .A(\_IFU_io_out_bits_instruction [20] ), .Z(\IDU/Control/_028_ ) );
BUF_X1 \IDU/Control/_244_ ( .A(\_IFU_io_out_bits_instruction [23] ), .Z(\IDU/Control/_031_ ) );
BUF_X1 \IDU/Control/_245_ ( .A(\_IFU_io_out_bits_instruction [22] ), .Z(\IDU/Control/_030_ ) );
BUF_X1 \IDU/Control/_246_ ( .A(\_IFU_io_out_bits_instruction [25] ), .Z(\IDU/Control/_033_ ) );
BUF_X1 \IDU/Control/_247_ ( .A(\_IFU_io_out_bits_instruction [24] ), .Z(\IDU/Control/_032_ ) );
BUF_X1 \IDU/Control/_248_ ( .A(\_IFU_io_out_bits_instruction [27] ), .Z(\IDU/Control/_035_ ) );
BUF_X1 \IDU/Control/_249_ ( .A(\_IFU_io_out_bits_instruction [26] ), .Z(\IDU/Control/_034_ ) );
BUF_X1 \IDU/Control/_250_ ( .A(\_IFU_io_out_bits_instruction [31] ), .Z(\IDU/Control/_040_ ) );
BUF_X1 \IDU/Control/_251_ ( .A(\IDU/Control/_009_ ), .Z(\_IDU_io_out_bits_control_csrCtr [0] ) );
BUF_X1 \IDU/Control/_252_ ( .A(\IDU/Control/_010_ ), .Z(\_IDU_io_out_bits_control_csrCtr [1] ) );
BUF_X1 \IDU/Control/_253_ ( .A(\IDU/Control/_011_ ), .Z(\_IDU_io_out_bits_control_csrCtr [2] ) );
BUF_X1 \IDU/Control/_254_ ( .A(\IDU/Control/_006_ ), .Z(\_IDU_io_out_bits_control_brType [0] ) );
BUF_X1 \IDU/Control/_255_ ( .A(\IDU/Control/_007_ ), .Z(\_IDU_io_out_bits_control_brType [1] ) );
BUF_X1 \IDU/Control/_256_ ( .A(\IDU/Control/_008_ ), .Z(\_IDU_io_out_bits_control_brType [2] ) );
BUF_X1 \IDU/Control/_257_ ( .A(\IDU/Control/_051_ ), .Z(_IDU_io_out_bits_control_pcSrc ) );
BUF_X1 \IDU/Control/_258_ ( .A(\IDU/Control/_049_ ), .Z(_IDU_io_out_bits_control_memRen ) );
BUF_X1 \IDU/Control/_259_ ( .A(\IDU/Control/_053_ ), .Z(\_IDU_io_out_bits_control_wbSrc [1] ) );
BUF_X1 \IDU/Control/_260_ ( .A(\IDU/Control/_048_ ), .Z(\IDU/_Control_io_isEnd ) );
BUF_X1 \IDU/Control/_261_ ( .A(\IDU/Control/_013_ ), .Z(\IDU/_Control_io_immType [0] ) );
BUF_X1 \IDU/Control/_262_ ( .A(\IDU/Control/_050_ ), .Z(_IDU_io_out_bits_control_memWen ) );
BUF_X1 \IDU/Control/_263_ ( .A(\IDU/Control/_014_ ), .Z(\IDU/_Control_io_immType [1] ) );
BUF_X1 \IDU/Control/_264_ ( .A(\IDU/Control/_015_ ), .Z(\IDU/_Control_io_immType [2] ) );
BUF_X1 \IDU/Control/_265_ ( .A(\IDU/Control/_002_ ), .Z(\_IDU_io_out_bits_control_aluBSrc [1] ) );
BUF_X1 \IDU/Control/_266_ ( .A(\IDU/Control/_052_ ), .Z(_IDU_io_out_bits_control_regWe ) );
BUF_X1 \IDU/Control/_267_ ( .A(\IDU/Control/_000_ ), .Z(_IDU_io_out_bits_control_aluASrc ) );
BUF_X1 \IDU/Control/_268_ ( .A(\IDU/Control/_001_ ), .Z(\_IDU_io_out_bits_control_aluBSrc [0] ) );
NOR2_X1 \IDU/ImmGen/_090_ ( .A1(\IDU/ImmGen/_000_ ), .A2(\IDU/ImmGen/_001_ ), .ZN(\IDU/ImmGen/_062_ ) );
INV_X32 \IDU/ImmGen/_091_ ( .A(\IDU/ImmGen/_002_ ), .ZN(\IDU/ImmGen/_063_ ) );
BUF_X4 \IDU/ImmGen/_092_ ( .A(\IDU/ImmGen/_063_ ), .Z(\IDU/ImmGen/_064_ ) );
NAND3_X1 \IDU/ImmGen/_093_ ( .A1(\IDU/ImmGen/_062_ ), .A2(\IDU/ImmGen/_064_ ), .A3(\IDU/ImmGen/_044_ ), .ZN(\IDU/ImmGen/_065_ ) );
INV_X4 \IDU/ImmGen/_094_ ( .A(\IDU/ImmGen/_000_ ), .ZN(\IDU/ImmGen/_066_ ) );
NAND4_X1 \IDU/ImmGen/_095_ ( .A1(\IDU/ImmGen/_064_ ), .A2(\IDU/ImmGen/_066_ ), .A3(\IDU/ImmGen/_001_ ), .A4(\IDU/ImmGen/_056_ ), .ZN(\IDU/ImmGen/_067_ ) );
NAND2_X1 \IDU/ImmGen/_096_ ( .A1(\IDU/ImmGen/_065_ ), .A2(\IDU/ImmGen/_067_ ), .ZN(\IDU/ImmGen/_003_ ) );
NAND3_X1 \IDU/ImmGen/_097_ ( .A1(\IDU/ImmGen/_064_ ), .A2(\IDU/ImmGen/_001_ ), .A3(\IDU/ImmGen/_057_ ), .ZN(\IDU/ImmGen/_068_ ) );
INV_X1 \IDU/ImmGen/_098_ ( .A(\IDU/ImmGen/_062_ ), .ZN(\IDU/ImmGen/_069_ ) );
INV_X1 \IDU/ImmGen/_099_ ( .A(\IDU/ImmGen/_045_ ), .ZN(\IDU/ImmGen/_070_ ) );
OAI21_X1 \IDU/ImmGen/_100_ ( .A(\IDU/ImmGen/_068_ ), .B1(\IDU/ImmGen/_069_ ), .B2(\IDU/ImmGen/_070_ ), .ZN(\IDU/ImmGen/_014_ ) );
NAND3_X1 \IDU/ImmGen/_101_ ( .A1(\IDU/ImmGen/_064_ ), .A2(\IDU/ImmGen/_001_ ), .A3(\IDU/ImmGen/_058_ ), .ZN(\IDU/ImmGen/_071_ ) );
INV_X1 \IDU/ImmGen/_102_ ( .A(\IDU/ImmGen/_046_ ), .ZN(\IDU/ImmGen/_072_ ) );
OAI21_X1 \IDU/ImmGen/_103_ ( .A(\IDU/ImmGen/_071_ ), .B1(\IDU/ImmGen/_069_ ), .B2(\IDU/ImmGen/_072_ ), .ZN(\IDU/ImmGen/_025_ ) );
NAND3_X1 \IDU/ImmGen/_104_ ( .A1(\IDU/ImmGen/_063_ ), .A2(\IDU/ImmGen/_001_ ), .A3(\IDU/ImmGen/_034_ ), .ZN(\IDU/ImmGen/_073_ ) );
INV_X1 \IDU/ImmGen/_105_ ( .A(\IDU/ImmGen/_047_ ), .ZN(\IDU/ImmGen/_074_ ) );
OAI21_X1 \IDU/ImmGen/_106_ ( .A(\IDU/ImmGen/_073_ ), .B1(\IDU/ImmGen/_069_ ), .B2(\IDU/ImmGen/_074_ ), .ZN(\IDU/ImmGen/_027_ ) );
NAND3_X1 \IDU/ImmGen/_107_ ( .A1(\IDU/ImmGen/_063_ ), .A2(\IDU/ImmGen/_001_ ), .A3(\IDU/ImmGen/_035_ ), .ZN(\IDU/ImmGen/_075_ ) );
INV_X1 \IDU/ImmGen/_108_ ( .A(\IDU/ImmGen/_048_ ), .ZN(\IDU/ImmGen/_076_ ) );
OAI21_X1 \IDU/ImmGen/_109_ ( .A(\IDU/ImmGen/_075_ ), .B1(\IDU/ImmGen/_069_ ), .B2(\IDU/ImmGen/_076_ ), .ZN(\IDU/ImmGen/_028_ ) );
INV_X1 \IDU/ImmGen/_110_ ( .A(\IDU/ImmGen/_049_ ), .ZN(\IDU/ImmGen/_077_ ) );
NOR2_X4 \IDU/ImmGen/_111_ ( .A1(\IDU/ImmGen/_066_ ), .A2(\IDU/ImmGen/_001_ ), .ZN(\IDU/ImmGen/_078_ ) );
AOI21_X1 \IDU/ImmGen/_112_ ( .A(\IDU/ImmGen/_077_ ), .B1(\IDU/ImmGen/_078_ ), .B2(\IDU/ImmGen/_064_ ), .ZN(\IDU/ImmGen/_029_ ) );
INV_X1 \IDU/ImmGen/_113_ ( .A(\IDU/ImmGen/_050_ ), .ZN(\IDU/ImmGen/_079_ ) );
AOI21_X1 \IDU/ImmGen/_114_ ( .A(\IDU/ImmGen/_079_ ), .B1(\IDU/ImmGen/_078_ ), .B2(\IDU/ImmGen/_064_ ), .ZN(\IDU/ImmGen/_030_ ) );
INV_X1 \IDU/ImmGen/_115_ ( .A(\IDU/ImmGen/_051_ ), .ZN(\IDU/ImmGen/_080_ ) );
AOI21_X1 \IDU/ImmGen/_116_ ( .A(\IDU/ImmGen/_080_ ), .B1(\IDU/ImmGen/_078_ ), .B2(\IDU/ImmGen/_064_ ), .ZN(\IDU/ImmGen/_031_ ) );
INV_X1 \IDU/ImmGen/_117_ ( .A(\IDU/ImmGen/_052_ ), .ZN(\IDU/ImmGen/_081_ ) );
AOI21_X1 \IDU/ImmGen/_118_ ( .A(\IDU/ImmGen/_081_ ), .B1(\IDU/ImmGen/_078_ ), .B2(\IDU/ImmGen/_064_ ), .ZN(\IDU/ImmGen/_032_ ) );
INV_X1 \IDU/ImmGen/_119_ ( .A(\IDU/ImmGen/_053_ ), .ZN(\IDU/ImmGen/_082_ ) );
AOI21_X1 \IDU/ImmGen/_120_ ( .A(\IDU/ImmGen/_082_ ), .B1(\IDU/ImmGen/_078_ ), .B2(\IDU/ImmGen/_064_ ), .ZN(\IDU/ImmGen/_033_ ) );
INV_X1 \IDU/ImmGen/_121_ ( .A(\IDU/ImmGen/_054_ ), .ZN(\IDU/ImmGen/_083_ ) );
AOI21_X1 \IDU/ImmGen/_122_ ( .A(\IDU/ImmGen/_083_ ), .B1(\IDU/ImmGen/_078_ ), .B2(\IDU/ImmGen/_064_ ), .ZN(\IDU/ImmGen/_004_ ) );
NAND4_X1 \IDU/ImmGen/_123_ ( .A1(\IDU/ImmGen/_063_ ), .A2(\IDU/ImmGen/_000_ ), .A3(\IDU/ImmGen/_001_ ), .A4(\IDU/ImmGen/_056_ ), .ZN(\IDU/ImmGen/_084_ ) );
AND2_X4 \IDU/ImmGen/_124_ ( .A1(\IDU/ImmGen/_078_ ), .A2(\IDU/ImmGen/_063_ ), .ZN(\IDU/ImmGen/_085_ ) );
NOR3_X4 \IDU/ImmGen/_125_ ( .A1(\IDU/ImmGen/_063_ ), .A2(\IDU/ImmGen/_000_ ), .A3(\IDU/ImmGen/_001_ ), .ZN(\IDU/ImmGen/_086_ ) );
NOR2_X4 \IDU/ImmGen/_126_ ( .A1(\IDU/ImmGen/_085_ ), .A2(\IDU/ImmGen/_086_ ), .ZN(\IDU/ImmGen/_087_ ) );
AOI22_X1 \IDU/ImmGen/_127_ ( .A1(\IDU/ImmGen/_087_ ), .A2(\IDU/ImmGen/_055_ ), .B1(\IDU/ImmGen/_044_ ), .B2(\IDU/ImmGen/_086_ ), .ZN(\IDU/ImmGen/_088_ ) );
AND3_X1 \IDU/ImmGen/_128_ ( .A1(\IDU/ImmGen/_063_ ), .A2(\IDU/ImmGen/_000_ ), .A3(\IDU/ImmGen/_001_ ), .ZN(\IDU/ImmGen/_089_ ) );
OAI21_X1 \IDU/ImmGen/_129_ ( .A(\IDU/ImmGen/_084_ ), .B1(\IDU/ImmGen/_088_ ), .B2(\IDU/ImmGen/_089_ ), .ZN(\IDU/ImmGen/_005_ ) );
MUX2_X1 \IDU/ImmGen/_130_ ( .A(\IDU/ImmGen/_036_ ), .B(\IDU/ImmGen/_055_ ), .S(\IDU/ImmGen/_087_ ), .Z(\IDU/ImmGen/_006_ ) );
MUX2_X1 \IDU/ImmGen/_131_ ( .A(\IDU/ImmGen/_037_ ), .B(\IDU/ImmGen/_055_ ), .S(\IDU/ImmGen/_087_ ), .Z(\IDU/ImmGen/_007_ ) );
MUX2_X1 \IDU/ImmGen/_132_ ( .A(\IDU/ImmGen/_038_ ), .B(\IDU/ImmGen/_055_ ), .S(\IDU/ImmGen/_087_ ), .Z(\IDU/ImmGen/_008_ ) );
MUX2_X1 \IDU/ImmGen/_133_ ( .A(\IDU/ImmGen/_039_ ), .B(\IDU/ImmGen/_055_ ), .S(\IDU/ImmGen/_087_ ), .Z(\IDU/ImmGen/_009_ ) );
MUX2_X1 \IDU/ImmGen/_134_ ( .A(\IDU/ImmGen/_040_ ), .B(\IDU/ImmGen/_055_ ), .S(\IDU/ImmGen/_087_ ), .Z(\IDU/ImmGen/_010_ ) );
MUX2_X1 \IDU/ImmGen/_135_ ( .A(\IDU/ImmGen/_041_ ), .B(\IDU/ImmGen/_055_ ), .S(\IDU/ImmGen/_087_ ), .Z(\IDU/ImmGen/_011_ ) );
MUX2_X1 \IDU/ImmGen/_136_ ( .A(\IDU/ImmGen/_042_ ), .B(\IDU/ImmGen/_055_ ), .S(\IDU/ImmGen/_087_ ), .Z(\IDU/ImmGen/_012_ ) );
MUX2_X1 \IDU/ImmGen/_137_ ( .A(\IDU/ImmGen/_043_ ), .B(\IDU/ImmGen/_055_ ), .S(\IDU/ImmGen/_087_ ), .Z(\IDU/ImmGen/_013_ ) );
MUX2_X1 \IDU/ImmGen/_138_ ( .A(\IDU/ImmGen/_055_ ), .B(\IDU/ImmGen/_044_ ), .S(\IDU/ImmGen/_085_ ), .Z(\IDU/ImmGen/_015_ ) );
INV_X1 \IDU/ImmGen/_139_ ( .A(\IDU/ImmGen/_085_ ), .ZN(\IDU/ImmGen/_059_ ) );
NAND2_X2 \IDU/ImmGen/_140_ ( .A1(\IDU/ImmGen/_059_ ), .A2(\IDU/ImmGen/_055_ ), .ZN(\IDU/ImmGen/_060_ ) );
BUF_X4 \IDU/ImmGen/_141_ ( .A(\IDU/ImmGen/_059_ ), .Z(\IDU/ImmGen/_061_ ) );
OAI21_X1 \IDU/ImmGen/_142_ ( .A(\IDU/ImmGen/_060_ ), .B1(\IDU/ImmGen/_070_ ), .B2(\IDU/ImmGen/_061_ ), .ZN(\IDU/ImmGen/_016_ ) );
OAI21_X1 \IDU/ImmGen/_143_ ( .A(\IDU/ImmGen/_060_ ), .B1(\IDU/ImmGen/_072_ ), .B2(\IDU/ImmGen/_061_ ), .ZN(\IDU/ImmGen/_017_ ) );
OAI21_X1 \IDU/ImmGen/_144_ ( .A(\IDU/ImmGen/_060_ ), .B1(\IDU/ImmGen/_074_ ), .B2(\IDU/ImmGen/_061_ ), .ZN(\IDU/ImmGen/_018_ ) );
OAI21_X1 \IDU/ImmGen/_145_ ( .A(\IDU/ImmGen/_060_ ), .B1(\IDU/ImmGen/_076_ ), .B2(\IDU/ImmGen/_061_ ), .ZN(\IDU/ImmGen/_019_ ) );
OAI21_X1 \IDU/ImmGen/_146_ ( .A(\IDU/ImmGen/_060_ ), .B1(\IDU/ImmGen/_077_ ), .B2(\IDU/ImmGen/_061_ ), .ZN(\IDU/ImmGen/_020_ ) );
OAI21_X1 \IDU/ImmGen/_147_ ( .A(\IDU/ImmGen/_060_ ), .B1(\IDU/ImmGen/_079_ ), .B2(\IDU/ImmGen/_061_ ), .ZN(\IDU/ImmGen/_021_ ) );
OAI21_X1 \IDU/ImmGen/_148_ ( .A(\IDU/ImmGen/_060_ ), .B1(\IDU/ImmGen/_080_ ), .B2(\IDU/ImmGen/_061_ ), .ZN(\IDU/ImmGen/_022_ ) );
OAI21_X1 \IDU/ImmGen/_149_ ( .A(\IDU/ImmGen/_060_ ), .B1(\IDU/ImmGen/_081_ ), .B2(\IDU/ImmGen/_061_ ), .ZN(\IDU/ImmGen/_023_ ) );
OAI21_X1 \IDU/ImmGen/_150_ ( .A(\IDU/ImmGen/_060_ ), .B1(\IDU/ImmGen/_082_ ), .B2(\IDU/ImmGen/_061_ ), .ZN(\IDU/ImmGen/_024_ ) );
OAI21_X1 \IDU/ImmGen/_151_ ( .A(\IDU/ImmGen/_060_ ), .B1(\IDU/ImmGen/_083_ ), .B2(\IDU/ImmGen/_061_ ), .ZN(\IDU/ImmGen/_026_ ) );
BUF_X1 \IDU/ImmGen/_152_ ( .A(\_IFU_io_out_bits_instruction [31] ), .Z(\_IDU_io_out_bits_imm [31] ) );
BUF_X1 \IDU/ImmGen/_153_ ( .A(\IDU/_Control_io_immType [2] ), .Z(\IDU/ImmGen/_002_ ) );
BUF_X1 \IDU/ImmGen/_154_ ( .A(\IDU/_Control_io_immType [0] ), .Z(\IDU/ImmGen/_000_ ) );
BUF_X1 \IDU/ImmGen/_155_ ( .A(\IDU/_Control_io_immType [1] ), .Z(\IDU/ImmGen/_001_ ) );
BUF_X1 \IDU/ImmGen/_156_ ( .A(\_IFU_io_out_bits_instruction [7] ), .Z(\IDU/ImmGen/_056_ ) );
BUF_X1 \IDU/ImmGen/_157_ ( .A(\_IFU_io_out_bits_instruction [20] ), .Z(\IDU/ImmGen/_044_ ) );
BUF_X1 \IDU/ImmGen/_158_ ( .A(\IDU/ImmGen/_003_ ), .Z(\_IDU_io_out_bits_imm [0] ) );
BUF_X1 \IDU/ImmGen/_159_ ( .A(\_IFU_io_out_bits_instruction [8] ), .Z(\IDU/ImmGen/_057_ ) );
BUF_X1 \IDU/ImmGen/_160_ ( .A(\_IFU_io_out_bits_instruction [21] ), .Z(\IDU/ImmGen/_045_ ) );
BUF_X1 \IDU/ImmGen/_161_ ( .A(\IDU/ImmGen/_014_ ), .Z(\_IDU_io_out_bits_imm [1] ) );
BUF_X1 \IDU/ImmGen/_162_ ( .A(\_IFU_io_out_bits_instruction [9] ), .Z(\IDU/ImmGen/_058_ ) );
BUF_X1 \IDU/ImmGen/_163_ ( .A(\_IFU_io_out_bits_instruction [22] ), .Z(\IDU/ImmGen/_046_ ) );
BUF_X1 \IDU/ImmGen/_164_ ( .A(\IDU/ImmGen/_025_ ), .Z(\_IDU_io_out_bits_imm [2] ) );
BUF_X1 \IDU/ImmGen/_165_ ( .A(\_IFU_io_out_bits_instruction [10] ), .Z(\IDU/ImmGen/_034_ ) );
BUF_X1 \IDU/ImmGen/_166_ ( .A(\_IFU_io_out_bits_instruction [23] ), .Z(\IDU/ImmGen/_047_ ) );
BUF_X1 \IDU/ImmGen/_167_ ( .A(\IDU/ImmGen/_027_ ), .Z(\_IDU_io_out_bits_imm [3] ) );
BUF_X1 \IDU/ImmGen/_168_ ( .A(\_IFU_io_out_bits_instruction [11] ), .Z(\IDU/ImmGen/_035_ ) );
BUF_X1 \IDU/ImmGen/_169_ ( .A(\_IFU_io_out_bits_instruction [24] ), .Z(\IDU/ImmGen/_048_ ) );
BUF_X1 \IDU/ImmGen/_170_ ( .A(\IDU/ImmGen/_028_ ), .Z(\_IDU_io_out_bits_imm [4] ) );
BUF_X1 \IDU/ImmGen/_171_ ( .A(\_IFU_io_out_bits_instruction [25] ), .Z(\IDU/ImmGen/_049_ ) );
BUF_X1 \IDU/ImmGen/_172_ ( .A(\IDU/ImmGen/_029_ ), .Z(\_IDU_io_out_bits_imm [5] ) );
BUF_X1 \IDU/ImmGen/_173_ ( .A(\_IFU_io_out_bits_instruction [26] ), .Z(\IDU/ImmGen/_050_ ) );
BUF_X1 \IDU/ImmGen/_174_ ( .A(\IDU/ImmGen/_030_ ), .Z(\_IDU_io_out_bits_imm [6] ) );
BUF_X1 \IDU/ImmGen/_175_ ( .A(\_IFU_io_out_bits_instruction [27] ), .Z(\IDU/ImmGen/_051_ ) );
BUF_X1 \IDU/ImmGen/_176_ ( .A(\IDU/ImmGen/_031_ ), .Z(\_IDU_io_out_bits_imm [7] ) );
BUF_X1 \IDU/ImmGen/_177_ ( .A(\_IFU_io_out_bits_instruction [28] ), .Z(\IDU/ImmGen/_052_ ) );
BUF_X1 \IDU/ImmGen/_178_ ( .A(\IDU/ImmGen/_032_ ), .Z(\_IDU_io_out_bits_imm [8] ) );
BUF_X1 \IDU/ImmGen/_179_ ( .A(\_IFU_io_out_bits_instruction [29] ), .Z(\IDU/ImmGen/_053_ ) );
BUF_X1 \IDU/ImmGen/_180_ ( .A(\IDU/ImmGen/_033_ ), .Z(\_IDU_io_out_bits_imm [9] ) );
BUF_X1 \IDU/ImmGen/_181_ ( .A(\_IFU_io_out_bits_instruction [30] ), .Z(\IDU/ImmGen/_054_ ) );
BUF_X1 \IDU/ImmGen/_182_ ( .A(\IDU/ImmGen/_004_ ), .Z(\_IDU_io_out_bits_imm [10] ) );
BUF_X1 \IDU/ImmGen/_183_ ( .A(\_IFU_io_out_bits_instruction [31] ), .Z(\IDU/ImmGen/_055_ ) );
BUF_X1 \IDU/ImmGen/_184_ ( .A(\IDU/ImmGen/_005_ ), .Z(\_IDU_io_out_bits_imm [11] ) );
BUF_X1 \IDU/ImmGen/_185_ ( .A(\_IFU_io_out_bits_instruction [12] ), .Z(\IDU/ImmGen/_036_ ) );
BUF_X1 \IDU/ImmGen/_186_ ( .A(\IDU/ImmGen/_006_ ), .Z(\_IDU_io_out_bits_imm [12] ) );
BUF_X1 \IDU/ImmGen/_187_ ( .A(\_IFU_io_out_bits_instruction [13] ), .Z(\IDU/ImmGen/_037_ ) );
BUF_X1 \IDU/ImmGen/_188_ ( .A(\IDU/ImmGen/_007_ ), .Z(\_IDU_io_out_bits_imm [13] ) );
BUF_X1 \IDU/ImmGen/_189_ ( .A(\_IFU_io_out_bits_instruction [14] ), .Z(\IDU/ImmGen/_038_ ) );
BUF_X1 \IDU/ImmGen/_190_ ( .A(\IDU/ImmGen/_008_ ), .Z(\_IDU_io_out_bits_imm [14] ) );
BUF_X1 \IDU/ImmGen/_191_ ( .A(\_IFU_io_out_bits_instruction [15] ), .Z(\IDU/ImmGen/_039_ ) );
BUF_X1 \IDU/ImmGen/_192_ ( .A(\IDU/ImmGen/_009_ ), .Z(\_IDU_io_out_bits_imm [15] ) );
BUF_X1 \IDU/ImmGen/_193_ ( .A(\_IFU_io_out_bits_instruction [16] ), .Z(\IDU/ImmGen/_040_ ) );
BUF_X1 \IDU/ImmGen/_194_ ( .A(\IDU/ImmGen/_010_ ), .Z(\_IDU_io_out_bits_imm [16] ) );
BUF_X1 \IDU/ImmGen/_195_ ( .A(\_IFU_io_out_bits_instruction [17] ), .Z(\IDU/ImmGen/_041_ ) );
BUF_X1 \IDU/ImmGen/_196_ ( .A(\IDU/ImmGen/_011_ ), .Z(\_IDU_io_out_bits_imm [17] ) );
BUF_X1 \IDU/ImmGen/_197_ ( .A(\_IFU_io_out_bits_instruction [18] ), .Z(\IDU/ImmGen/_042_ ) );
BUF_X1 \IDU/ImmGen/_198_ ( .A(\IDU/ImmGen/_012_ ), .Z(\_IDU_io_out_bits_imm [18] ) );
BUF_X1 \IDU/ImmGen/_199_ ( .A(\_IFU_io_out_bits_instruction [19] ), .Z(\IDU/ImmGen/_043_ ) );
BUF_X1 \IDU/ImmGen/_200_ ( .A(\IDU/ImmGen/_013_ ), .Z(\_IDU_io_out_bits_imm [19] ) );
BUF_X1 \IDU/ImmGen/_201_ ( .A(\IDU/ImmGen/_015_ ), .Z(\_IDU_io_out_bits_imm [20] ) );
BUF_X1 \IDU/ImmGen/_202_ ( .A(\IDU/ImmGen/_016_ ), .Z(\_IDU_io_out_bits_imm [21] ) );
BUF_X1 \IDU/ImmGen/_203_ ( .A(\IDU/ImmGen/_017_ ), .Z(\_IDU_io_out_bits_imm [22] ) );
BUF_X1 \IDU/ImmGen/_204_ ( .A(\IDU/ImmGen/_018_ ), .Z(\_IDU_io_out_bits_imm [23] ) );
BUF_X1 \IDU/ImmGen/_205_ ( .A(\IDU/ImmGen/_019_ ), .Z(\_IDU_io_out_bits_imm [24] ) );
BUF_X1 \IDU/ImmGen/_206_ ( .A(\IDU/ImmGen/_020_ ), .Z(\_IDU_io_out_bits_imm [25] ) );
BUF_X1 \IDU/ImmGen/_207_ ( .A(\IDU/ImmGen/_021_ ), .Z(\_IDU_io_out_bits_imm [26] ) );
BUF_X1 \IDU/ImmGen/_208_ ( .A(\IDU/ImmGen/_022_ ), .Z(\_IDU_io_out_bits_imm [27] ) );
BUF_X1 \IDU/ImmGen/_209_ ( .A(\IDU/ImmGen/_023_ ), .Z(\_IDU_io_out_bits_imm [28] ) );
BUF_X1 \IDU/ImmGen/_210_ ( .A(\IDU/ImmGen/_024_ ), .Z(\_IDU_io_out_bits_imm [29] ) );
BUF_X1 \IDU/ImmGen/_211_ ( .A(\IDU/ImmGen/_026_ ), .Z(\_IDU_io_out_bits_imm [30] ) );
AND2_X1 \IFU/_424_ ( .A1(\IFU/_290_ ), .A2(\IFU/_291_ ), .ZN(\IFU/_201_ ) );
INV_X32 \IFU/_425_ ( .A(\IFU/_290_ ), .ZN(\IFU/_202_ ) );
AND2_X4 \IFU/_426_ ( .A1(\IFU/_202_ ), .A2(\IFU/_291_ ), .ZN(\IFU/_166_ ) );
NOR2_X1 \IFU/_427_ ( .A1(\IFU/_202_ ), .A2(\IFU/_291_ ), .ZN(\IFU/_133_ ) );
NOR2_X4 \IFU/_428_ ( .A1(\IFU/_290_ ), .A2(\IFU/_291_ ), .ZN(\IFU/_098_ ) );
AND2_X4 \IFU/_429_ ( .A1(\IFU/_166_ ), .A2(\IFU/_167_ ), .ZN(\IFU/_203_ ) );
BUF_X8 \IFU/_430_ ( .A(\IFU/_203_ ), .Z(\IFU/_204_ ) );
INV_X1 \IFU/_431_ ( .A(\IFU/_204_ ), .ZN(\IFU/_205_ ) );
INV_X1 \IFU/_432_ ( .A(\IFU/_289_ ), .ZN(\IFU/_206_ ) );
CLKBUF_X2 \IFU/_433_ ( .A(\IFU/_206_ ), .Z(\IFU/_207_ ) );
OR3_X1 \IFU/_434_ ( .A1(\IFU/_202_ ), .A2(\IFU/_291_ ), .A3(\IFU/_132_ ), .ZN(\IFU/_208_ ) );
INV_X1 \IFU/_435_ ( .A(\IFU/_200_ ), .ZN(\IFU/_209_ ) );
AOI22_X1 \IFU/_436_ ( .A1(\IFU/_209_ ), .A2(\IFU/_201_ ), .B1(\IFU/_098_ ), .B2(\IFU/_099_ ), .ZN(\IFU/_210_ ) );
NAND4_X1 \IFU/_437_ ( .A1(\IFU/_205_ ), .A2(\IFU/_207_ ), .A3(\IFU/_208_ ), .A4(\IFU/_210_ ), .ZN(\IFU/_000_ ) );
AOI221_X4 \IFU/_438_ ( .A(\IFU/_166_ ), .B1(\IFU/_201_ ), .B2(\IFU/_209_ ), .C1(\IFU/_132_ ), .C2(\IFU/_133_ ), .ZN(\IFU/_211_ ) );
NOR2_X1 \IFU/_439_ ( .A1(\IFU/_211_ ), .A2(\IFU/_289_ ), .ZN(\IFU/_001_ ) );
AND2_X4 \IFU/_440_ ( .A1(\IFU/_098_ ), .A2(\IFU/_099_ ), .ZN(\IFU/_212_ ) );
BUF_X8 \IFU/_441_ ( .A(\IFU/_212_ ), .Z(\IFU/_213_ ) );
MUX2_X1 \IFU/_442_ ( .A(\IFU/_100_ ), .B(\IFU/_066_ ), .S(\IFU/_213_ ), .Z(\IFU/_214_ ) );
AND2_X1 \IFU/_443_ ( .A1(\IFU/_214_ ), .A2(\IFU/_207_ ), .ZN(\IFU/_002_ ) );
MUX2_X1 \IFU/_444_ ( .A(\IFU/_111_ ), .B(\IFU/_077_ ), .S(\IFU/_213_ ), .Z(\IFU/_215_ ) );
AND2_X1 \IFU/_445_ ( .A1(\IFU/_215_ ), .A2(\IFU/_207_ ), .ZN(\IFU/_003_ ) );
MUX2_X1 \IFU/_446_ ( .A(\IFU/_122_ ), .B(\IFU/_088_ ), .S(\IFU/_213_ ), .Z(\IFU/_216_ ) );
AND2_X1 \IFU/_447_ ( .A1(\IFU/_216_ ), .A2(\IFU/_207_ ), .ZN(\IFU/_004_ ) );
MUX2_X1 \IFU/_448_ ( .A(\IFU/_125_ ), .B(\IFU/_091_ ), .S(\IFU/_213_ ), .Z(\IFU/_217_ ) );
AND2_X1 \IFU/_449_ ( .A1(\IFU/_217_ ), .A2(\IFU/_207_ ), .ZN(\IFU/_005_ ) );
MUX2_X1 \IFU/_450_ ( .A(\IFU/_126_ ), .B(\IFU/_092_ ), .S(\IFU/_213_ ), .Z(\IFU/_218_ ) );
AND2_X1 \IFU/_451_ ( .A1(\IFU/_218_ ), .A2(\IFU/_207_ ), .ZN(\IFU/_006_ ) );
MUX2_X1 \IFU/_452_ ( .A(\IFU/_127_ ), .B(\IFU/_093_ ), .S(\IFU/_213_ ), .Z(\IFU/_219_ ) );
AND2_X1 \IFU/_453_ ( .A1(\IFU/_219_ ), .A2(\IFU/_207_ ), .ZN(\IFU/_007_ ) );
MUX2_X1 \IFU/_454_ ( .A(\IFU/_128_ ), .B(\IFU/_094_ ), .S(\IFU/_213_ ), .Z(\IFU/_220_ ) );
AND2_X1 \IFU/_455_ ( .A1(\IFU/_220_ ), .A2(\IFU/_207_ ), .ZN(\IFU/_008_ ) );
MUX2_X1 \IFU/_456_ ( .A(\IFU/_129_ ), .B(\IFU/_095_ ), .S(\IFU/_213_ ), .Z(\IFU/_221_ ) );
AND2_X1 \IFU/_457_ ( .A1(\IFU/_221_ ), .A2(\IFU/_207_ ), .ZN(\IFU/_009_ ) );
MUX2_X1 \IFU/_458_ ( .A(\IFU/_130_ ), .B(\IFU/_096_ ), .S(\IFU/_213_ ), .Z(\IFU/_222_ ) );
CLKBUF_X2 \IFU/_459_ ( .A(\IFU/_206_ ), .Z(\IFU/_223_ ) );
AND2_X1 \IFU/_460_ ( .A1(\IFU/_222_ ), .A2(\IFU/_223_ ), .ZN(\IFU/_010_ ) );
MUX2_X1 \IFU/_461_ ( .A(\IFU/_131_ ), .B(\IFU/_097_ ), .S(\IFU/_213_ ), .Z(\IFU/_224_ ) );
AND2_X1 \IFU/_462_ ( .A1(\IFU/_224_ ), .A2(\IFU/_223_ ), .ZN(\IFU/_011_ ) );
BUF_X8 \IFU/_463_ ( .A(\IFU/_212_ ), .Z(\IFU/_225_ ) );
MUX2_X1 \IFU/_464_ ( .A(\IFU/_101_ ), .B(\IFU/_067_ ), .S(\IFU/_225_ ), .Z(\IFU/_226_ ) );
AND2_X1 \IFU/_465_ ( .A1(\IFU/_226_ ), .A2(\IFU/_223_ ), .ZN(\IFU/_012_ ) );
MUX2_X1 \IFU/_466_ ( .A(\IFU/_102_ ), .B(\IFU/_068_ ), .S(\IFU/_225_ ), .Z(\IFU/_227_ ) );
AND2_X1 \IFU/_467_ ( .A1(\IFU/_227_ ), .A2(\IFU/_223_ ), .ZN(\IFU/_013_ ) );
MUX2_X1 \IFU/_468_ ( .A(\IFU/_103_ ), .B(\IFU/_069_ ), .S(\IFU/_225_ ), .Z(\IFU/_228_ ) );
AND2_X1 \IFU/_469_ ( .A1(\IFU/_228_ ), .A2(\IFU/_223_ ), .ZN(\IFU/_014_ ) );
MUX2_X1 \IFU/_470_ ( .A(\IFU/_104_ ), .B(\IFU/_070_ ), .S(\IFU/_225_ ), .Z(\IFU/_229_ ) );
AND2_X1 \IFU/_471_ ( .A1(\IFU/_229_ ), .A2(\IFU/_223_ ), .ZN(\IFU/_015_ ) );
MUX2_X1 \IFU/_472_ ( .A(\IFU/_105_ ), .B(\IFU/_071_ ), .S(\IFU/_225_ ), .Z(\IFU/_230_ ) );
AND2_X1 \IFU/_473_ ( .A1(\IFU/_230_ ), .A2(\IFU/_223_ ), .ZN(\IFU/_016_ ) );
MUX2_X1 \IFU/_474_ ( .A(\IFU/_106_ ), .B(\IFU/_072_ ), .S(\IFU/_225_ ), .Z(\IFU/_231_ ) );
AND2_X1 \IFU/_475_ ( .A1(\IFU/_231_ ), .A2(\IFU/_223_ ), .ZN(\IFU/_017_ ) );
MUX2_X1 \IFU/_476_ ( .A(\IFU/_107_ ), .B(\IFU/_073_ ), .S(\IFU/_225_ ), .Z(\IFU/_232_ ) );
AND2_X1 \IFU/_477_ ( .A1(\IFU/_232_ ), .A2(\IFU/_223_ ), .ZN(\IFU/_018_ ) );
MUX2_X1 \IFU/_478_ ( .A(\IFU/_108_ ), .B(\IFU/_074_ ), .S(\IFU/_225_ ), .Z(\IFU/_233_ ) );
AND2_X1 \IFU/_479_ ( .A1(\IFU/_233_ ), .A2(\IFU/_223_ ), .ZN(\IFU/_019_ ) );
MUX2_X1 \IFU/_480_ ( .A(\IFU/_109_ ), .B(\IFU/_075_ ), .S(\IFU/_225_ ), .Z(\IFU/_234_ ) );
CLKBUF_X2 \IFU/_481_ ( .A(\IFU/_206_ ), .Z(\IFU/_235_ ) );
AND2_X1 \IFU/_482_ ( .A1(\IFU/_234_ ), .A2(\IFU/_235_ ), .ZN(\IFU/_020_ ) );
MUX2_X1 \IFU/_483_ ( .A(\IFU/_110_ ), .B(\IFU/_076_ ), .S(\IFU/_225_ ), .Z(\IFU/_236_ ) );
AND2_X1 \IFU/_484_ ( .A1(\IFU/_236_ ), .A2(\IFU/_235_ ), .ZN(\IFU/_021_ ) );
BUF_X8 \IFU/_485_ ( .A(\IFU/_212_ ), .Z(\IFU/_237_ ) );
MUX2_X1 \IFU/_486_ ( .A(\IFU/_112_ ), .B(\IFU/_078_ ), .S(\IFU/_237_ ), .Z(\IFU/_238_ ) );
AND2_X1 \IFU/_487_ ( .A1(\IFU/_238_ ), .A2(\IFU/_235_ ), .ZN(\IFU/_022_ ) );
MUX2_X1 \IFU/_488_ ( .A(\IFU/_113_ ), .B(\IFU/_079_ ), .S(\IFU/_237_ ), .Z(\IFU/_239_ ) );
AND2_X1 \IFU/_489_ ( .A1(\IFU/_239_ ), .A2(\IFU/_235_ ), .ZN(\IFU/_023_ ) );
MUX2_X1 \IFU/_490_ ( .A(\IFU/_114_ ), .B(\IFU/_080_ ), .S(\IFU/_237_ ), .Z(\IFU/_240_ ) );
AND2_X1 \IFU/_491_ ( .A1(\IFU/_240_ ), .A2(\IFU/_235_ ), .ZN(\IFU/_024_ ) );
MUX2_X1 \IFU/_492_ ( .A(\IFU/_115_ ), .B(\IFU/_081_ ), .S(\IFU/_237_ ), .Z(\IFU/_241_ ) );
AND2_X1 \IFU/_493_ ( .A1(\IFU/_241_ ), .A2(\IFU/_235_ ), .ZN(\IFU/_025_ ) );
MUX2_X1 \IFU/_494_ ( .A(\IFU/_116_ ), .B(\IFU/_082_ ), .S(\IFU/_237_ ), .Z(\IFU/_242_ ) );
AND2_X1 \IFU/_495_ ( .A1(\IFU/_242_ ), .A2(\IFU/_235_ ), .ZN(\IFU/_026_ ) );
MUX2_X1 \IFU/_496_ ( .A(\IFU/_117_ ), .B(\IFU/_083_ ), .S(\IFU/_237_ ), .Z(\IFU/_243_ ) );
AND2_X1 \IFU/_497_ ( .A1(\IFU/_243_ ), .A2(\IFU/_235_ ), .ZN(\IFU/_027_ ) );
MUX2_X1 \IFU/_498_ ( .A(\IFU/_118_ ), .B(\IFU/_084_ ), .S(\IFU/_237_ ), .Z(\IFU/_244_ ) );
AND2_X1 \IFU/_499_ ( .A1(\IFU/_244_ ), .A2(\IFU/_235_ ), .ZN(\IFU/_028_ ) );
MUX2_X1 \IFU/_500_ ( .A(\IFU/_119_ ), .B(\IFU/_085_ ), .S(\IFU/_237_ ), .Z(\IFU/_245_ ) );
AND2_X1 \IFU/_501_ ( .A1(\IFU/_245_ ), .A2(\IFU/_235_ ), .ZN(\IFU/_029_ ) );
MUX2_X1 \IFU/_502_ ( .A(\IFU/_120_ ), .B(\IFU/_086_ ), .S(\IFU/_212_ ), .Z(\IFU/_246_ ) );
OR2_X1 \IFU/_503_ ( .A1(\IFU/_246_ ), .A2(\IFU/_289_ ), .ZN(\IFU/_030_ ) );
MUX2_X1 \IFU/_504_ ( .A(\IFU/_121_ ), .B(\IFU/_087_ ), .S(\IFU/_212_ ), .Z(\IFU/_247_ ) );
OR2_X1 \IFU/_505_ ( .A1(\IFU/_247_ ), .A2(\IFU/_289_ ), .ZN(\IFU/_031_ ) );
MUX2_X1 \IFU/_506_ ( .A(\IFU/_123_ ), .B(\IFU/_089_ ), .S(\IFU/_237_ ), .Z(\IFU/_248_ ) );
CLKBUF_X2 \IFU/_507_ ( .A(\IFU/_206_ ), .Z(\IFU/_249_ ) );
AND2_X1 \IFU/_508_ ( .A1(\IFU/_248_ ), .A2(\IFU/_249_ ), .ZN(\IFU/_032_ ) );
MUX2_X1 \IFU/_509_ ( .A(\IFU/_124_ ), .B(\IFU/_090_ ), .S(\IFU/_237_ ), .Z(\IFU/_250_ ) );
AND2_X1 \IFU/_510_ ( .A1(\IFU/_250_ ), .A2(\IFU/_249_ ), .ZN(\IFU/_033_ ) );
OR2_X2 \IFU/_511_ ( .A1(\IFU/_205_ ), .A2(\IFU/_134_ ), .ZN(\IFU/_251_ ) );
BUF_X8 \IFU/_512_ ( .A(\IFU/_204_ ), .Z(\IFU/_252_ ) );
OAI211_X2 \IFU/_513_ ( .A(\IFU/_251_ ), .B(\IFU/_206_ ), .C1(\IFU/_168_ ), .C2(\IFU/_252_ ), .ZN(\IFU/_253_ ) );
NAND2_X1 \IFU/_514_ ( .A1(\IFU/_253_ ), .A2(\IFU/_207_ ), .ZN(\IFU/_034_ ) );
MUX2_X1 \IFU/_515_ ( .A(\IFU/_179_ ), .B(\IFU/_145_ ), .S(\IFU/_204_ ), .Z(\IFU/_254_ ) );
OR2_X1 \IFU/_516_ ( .A1(\IFU/_254_ ), .A2(\IFU/_289_ ), .ZN(\IFU/_035_ ) );
MUX2_X1 \IFU/_517_ ( .A(\IFU/_190_ ), .B(\IFU/_156_ ), .S(\IFU/_252_ ), .Z(\IFU/_255_ ) );
AND2_X1 \IFU/_518_ ( .A1(\IFU/_255_ ), .A2(\IFU/_249_ ), .ZN(\IFU/_036_ ) );
MUX2_X1 \IFU/_519_ ( .A(\IFU/_193_ ), .B(\IFU/_159_ ), .S(\IFU/_252_ ), .Z(\IFU/_256_ ) );
AND2_X1 \IFU/_520_ ( .A1(\IFU/_256_ ), .A2(\IFU/_249_ ), .ZN(\IFU/_037_ ) );
MUX2_X1 \IFU/_521_ ( .A(\IFU/_194_ ), .B(\IFU/_160_ ), .S(\IFU/_204_ ), .Z(\IFU/_257_ ) );
OR2_X1 \IFU/_522_ ( .A1(\IFU/_257_ ), .A2(\IFU/_289_ ), .ZN(\IFU/_038_ ) );
MUX2_X1 \IFU/_523_ ( .A(\IFU/_195_ ), .B(\IFU/_161_ ), .S(\IFU/_252_ ), .Z(\IFU/_258_ ) );
AND2_X1 \IFU/_524_ ( .A1(\IFU/_258_ ), .A2(\IFU/_249_ ), .ZN(\IFU/_039_ ) );
MUX2_X1 \IFU/_525_ ( .A(\IFU/_196_ ), .B(\IFU/_162_ ), .S(\IFU/_252_ ), .Z(\IFU/_259_ ) );
AND2_X1 \IFU/_526_ ( .A1(\IFU/_259_ ), .A2(\IFU/_249_ ), .ZN(\IFU/_040_ ) );
MUX2_X1 \IFU/_527_ ( .A(\IFU/_197_ ), .B(\IFU/_163_ ), .S(\IFU/_252_ ), .Z(\IFU/_260_ ) );
AND2_X1 \IFU/_528_ ( .A1(\IFU/_260_ ), .A2(\IFU/_249_ ), .ZN(\IFU/_041_ ) );
MUX2_X1 \IFU/_529_ ( .A(\IFU/_198_ ), .B(\IFU/_164_ ), .S(\IFU/_252_ ), .Z(\IFU/_261_ ) );
AND2_X1 \IFU/_530_ ( .A1(\IFU/_261_ ), .A2(\IFU/_249_ ), .ZN(\IFU/_042_ ) );
MUX2_X1 \IFU/_531_ ( .A(\IFU/_199_ ), .B(\IFU/_165_ ), .S(\IFU/_252_ ), .Z(\IFU/_262_ ) );
AND2_X1 \IFU/_532_ ( .A1(\IFU/_262_ ), .A2(\IFU/_249_ ), .ZN(\IFU/_043_ ) );
MUX2_X1 \IFU/_533_ ( .A(\IFU/_169_ ), .B(\IFU/_135_ ), .S(\IFU/_252_ ), .Z(\IFU/_263_ ) );
AND2_X1 \IFU/_534_ ( .A1(\IFU/_263_ ), .A2(\IFU/_249_ ), .ZN(\IFU/_044_ ) );
MUX2_X1 \IFU/_535_ ( .A(\IFU/_170_ ), .B(\IFU/_136_ ), .S(\IFU/_252_ ), .Z(\IFU/_264_ ) );
CLKBUF_X2 \IFU/_536_ ( .A(\IFU/_206_ ), .Z(\IFU/_265_ ) );
AND2_X1 \IFU/_537_ ( .A1(\IFU/_264_ ), .A2(\IFU/_265_ ), .ZN(\IFU/_045_ ) );
BUF_X8 \IFU/_538_ ( .A(\IFU/_204_ ), .Z(\IFU/_266_ ) );
MUX2_X1 \IFU/_539_ ( .A(\IFU/_171_ ), .B(\IFU/_137_ ), .S(\IFU/_266_ ), .Z(\IFU/_267_ ) );
AND2_X1 \IFU/_540_ ( .A1(\IFU/_267_ ), .A2(\IFU/_265_ ), .ZN(\IFU/_046_ ) );
MUX2_X1 \IFU/_541_ ( .A(\IFU/_172_ ), .B(\IFU/_138_ ), .S(\IFU/_266_ ), .Z(\IFU/_268_ ) );
AND2_X1 \IFU/_542_ ( .A1(\IFU/_268_ ), .A2(\IFU/_265_ ), .ZN(\IFU/_047_ ) );
MUX2_X1 \IFU/_543_ ( .A(\IFU/_173_ ), .B(\IFU/_139_ ), .S(\IFU/_266_ ), .Z(\IFU/_269_ ) );
AND2_X1 \IFU/_544_ ( .A1(\IFU/_269_ ), .A2(\IFU/_265_ ), .ZN(\IFU/_048_ ) );
MUX2_X1 \IFU/_545_ ( .A(\IFU/_174_ ), .B(\IFU/_140_ ), .S(\IFU/_266_ ), .Z(\IFU/_270_ ) );
AND2_X1 \IFU/_546_ ( .A1(\IFU/_270_ ), .A2(\IFU/_265_ ), .ZN(\IFU/_049_ ) );
MUX2_X1 \IFU/_547_ ( .A(\IFU/_175_ ), .B(\IFU/_141_ ), .S(\IFU/_266_ ), .Z(\IFU/_271_ ) );
AND2_X1 \IFU/_548_ ( .A1(\IFU/_271_ ), .A2(\IFU/_265_ ), .ZN(\IFU/_050_ ) );
MUX2_X1 \IFU/_549_ ( .A(\IFU/_176_ ), .B(\IFU/_142_ ), .S(\IFU/_266_ ), .Z(\IFU/_272_ ) );
AND2_X1 \IFU/_550_ ( .A1(\IFU/_272_ ), .A2(\IFU/_265_ ), .ZN(\IFU/_051_ ) );
MUX2_X1 \IFU/_551_ ( .A(\IFU/_177_ ), .B(\IFU/_143_ ), .S(\IFU/_266_ ), .Z(\IFU/_273_ ) );
AND2_X1 \IFU/_552_ ( .A1(\IFU/_273_ ), .A2(\IFU/_265_ ), .ZN(\IFU/_052_ ) );
MUX2_X1 \IFU/_553_ ( .A(\IFU/_178_ ), .B(\IFU/_144_ ), .S(\IFU/_266_ ), .Z(\IFU/_274_ ) );
AND2_X1 \IFU/_554_ ( .A1(\IFU/_274_ ), .A2(\IFU/_265_ ), .ZN(\IFU/_053_ ) );
MUX2_X1 \IFU/_555_ ( .A(\IFU/_180_ ), .B(\IFU/_146_ ), .S(\IFU/_266_ ), .Z(\IFU/_275_ ) );
AND2_X1 \IFU/_556_ ( .A1(\IFU/_275_ ), .A2(\IFU/_265_ ), .ZN(\IFU/_054_ ) );
MUX2_X1 \IFU/_557_ ( .A(\IFU/_181_ ), .B(\IFU/_147_ ), .S(\IFU/_266_ ), .Z(\IFU/_276_ ) );
CLKBUF_X2 \IFU/_558_ ( .A(\IFU/_206_ ), .Z(\IFU/_277_ ) );
AND2_X1 \IFU/_559_ ( .A1(\IFU/_276_ ), .A2(\IFU/_277_ ), .ZN(\IFU/_055_ ) );
BUF_X8 \IFU/_560_ ( .A(\IFU/_204_ ), .Z(\IFU/_278_ ) );
MUX2_X1 \IFU/_561_ ( .A(\IFU/_182_ ), .B(\IFU/_148_ ), .S(\IFU/_278_ ), .Z(\IFU/_279_ ) );
AND2_X1 \IFU/_562_ ( .A1(\IFU/_279_ ), .A2(\IFU/_277_ ), .ZN(\IFU/_056_ ) );
MUX2_X1 \IFU/_563_ ( .A(\IFU/_183_ ), .B(\IFU/_149_ ), .S(\IFU/_278_ ), .Z(\IFU/_280_ ) );
AND2_X1 \IFU/_564_ ( .A1(\IFU/_280_ ), .A2(\IFU/_277_ ), .ZN(\IFU/_057_ ) );
MUX2_X1 \IFU/_565_ ( .A(\IFU/_184_ ), .B(\IFU/_150_ ), .S(\IFU/_278_ ), .Z(\IFU/_281_ ) );
AND2_X1 \IFU/_566_ ( .A1(\IFU/_281_ ), .A2(\IFU/_277_ ), .ZN(\IFU/_058_ ) );
MUX2_X1 \IFU/_567_ ( .A(\IFU/_185_ ), .B(\IFU/_151_ ), .S(\IFU/_278_ ), .Z(\IFU/_282_ ) );
AND2_X1 \IFU/_568_ ( .A1(\IFU/_282_ ), .A2(\IFU/_277_ ), .ZN(\IFU/_059_ ) );
MUX2_X1 \IFU/_569_ ( .A(\IFU/_186_ ), .B(\IFU/_152_ ), .S(\IFU/_278_ ), .Z(\IFU/_283_ ) );
AND2_X1 \IFU/_570_ ( .A1(\IFU/_283_ ), .A2(\IFU/_277_ ), .ZN(\IFU/_060_ ) );
MUX2_X1 \IFU/_571_ ( .A(\IFU/_187_ ), .B(\IFU/_153_ ), .S(\IFU/_278_ ), .Z(\IFU/_284_ ) );
AND2_X1 \IFU/_572_ ( .A1(\IFU/_284_ ), .A2(\IFU/_277_ ), .ZN(\IFU/_061_ ) );
MUX2_X1 \IFU/_573_ ( .A(\IFU/_188_ ), .B(\IFU/_154_ ), .S(\IFU/_278_ ), .Z(\IFU/_285_ ) );
AND2_X1 \IFU/_574_ ( .A1(\IFU/_285_ ), .A2(\IFU/_277_ ), .ZN(\IFU/_062_ ) );
MUX2_X1 \IFU/_575_ ( .A(\IFU/_189_ ), .B(\IFU/_155_ ), .S(\IFU/_278_ ), .Z(\IFU/_286_ ) );
AND2_X1 \IFU/_576_ ( .A1(\IFU/_286_ ), .A2(\IFU/_277_ ), .ZN(\IFU/_063_ ) );
MUX2_X1 \IFU/_577_ ( .A(\IFU/_191_ ), .B(\IFU/_157_ ), .S(\IFU/_278_ ), .Z(\IFU/_287_ ) );
AND2_X1 \IFU/_578_ ( .A1(\IFU/_287_ ), .A2(\IFU/_277_ ), .ZN(\IFU/_064_ ) );
MUX2_X1 \IFU/_579_ ( .A(\IFU/_192_ ), .B(\IFU/_158_ ), .S(\IFU/_278_ ), .Z(\IFU/_288_ ) );
AND2_X1 \IFU/_580_ ( .A1(\IFU/_288_ ), .A2(\IFU/_206_ ), .ZN(\IFU/_065_ ) );
DFF_X1 \IFU/_581_ ( .D(\IFU/_358_ ), .CK(clock ), .Q(\IFU/state [0] ), .QN(\IFU/_357_ ) );
DFF_X1 \IFU/_582_ ( .D(\IFU/_359_ ), .CK(clock ), .Q(\IFU/state [1] ), .QN(\IFU/_356_ ) );
DFF_X1 \IFU/_583_ ( .D(\IFU/_360_ ), .CK(clock ), .Q(\_IFU_io_master_araddr [0] ), .QN(\IFU/_355_ ) );
DFF_X1 \IFU/_584_ ( .D(\IFU/_361_ ), .CK(clock ), .Q(\_IFU_io_master_araddr [1] ), .QN(\IFU/_354_ ) );
DFF_X1 \IFU/_585_ ( .D(\IFU/_362_ ), .CK(clock ), .Q(\_IFU_io_master_araddr [2] ), .QN(\IFU/_353_ ) );
DFF_X1 \IFU/_586_ ( .D(\IFU/_363_ ), .CK(clock ), .Q(\_IFU_io_master_araddr [3] ), .QN(\IFU/_352_ ) );
DFF_X1 \IFU/_587_ ( .D(\IFU/_364_ ), .CK(clock ), .Q(\_IFU_io_master_araddr [4] ), .QN(\IFU/_351_ ) );
DFF_X1 \IFU/_588_ ( .D(\IFU/_365_ ), .CK(clock ), .Q(\_IFU_io_master_araddr [5] ), .QN(\IFU/_350_ ) );
DFF_X1 \IFU/_589_ ( .D(\IFU/_366_ ), .CK(clock ), .Q(\_IFU_io_master_araddr [6] ), .QN(\IFU/_349_ ) );
DFF_X1 \IFU/_590_ ( .D(\IFU/_367_ ), .CK(clock ), .Q(\_IFU_io_master_araddr [7] ), .QN(\IFU/_348_ ) );
DFF_X1 \IFU/_591_ ( .D(\IFU/_368_ ), .CK(clock ), .Q(\_IFU_io_master_araddr [8] ), .QN(\IFU/_347_ ) );
DFF_X1 \IFU/_592_ ( .D(\IFU/_369_ ), .CK(clock ), .Q(\_IFU_io_master_araddr [9] ), .QN(\IFU/_346_ ) );
DFF_X1 \IFU/_593_ ( .D(\IFU/_370_ ), .CK(clock ), .Q(\_IFU_io_master_araddr [10] ), .QN(\IFU/_345_ ) );
DFF_X1 \IFU/_594_ ( .D(\IFU/_371_ ), .CK(clock ), .Q(\_IFU_io_master_araddr [11] ), .QN(\IFU/_344_ ) );
DFF_X1 \IFU/_595_ ( .D(\IFU/_372_ ), .CK(clock ), .Q(\_IFU_io_master_araddr [12] ), .QN(\IFU/_343_ ) );
DFF_X1 \IFU/_596_ ( .D(\IFU/_373_ ), .CK(clock ), .Q(\_IFU_io_master_araddr [13] ), .QN(\IFU/_342_ ) );
DFF_X1 \IFU/_597_ ( .D(\IFU/_374_ ), .CK(clock ), .Q(\_IFU_io_master_araddr [14] ), .QN(\IFU/_341_ ) );
DFF_X1 \IFU/_598_ ( .D(\IFU/_375_ ), .CK(clock ), .Q(\_IFU_io_master_araddr [15] ), .QN(\IFU/_340_ ) );
DFF_X1 \IFU/_599_ ( .D(\IFU/_376_ ), .CK(clock ), .Q(\_IFU_io_master_araddr [16] ), .QN(\IFU/_339_ ) );
DFF_X1 \IFU/_600_ ( .D(\IFU/_377_ ), .CK(clock ), .Q(\_IFU_io_master_araddr [17] ), .QN(\IFU/_338_ ) );
DFF_X1 \IFU/_601_ ( .D(\IFU/_378_ ), .CK(clock ), .Q(\_IFU_io_master_araddr [18] ), .QN(\IFU/_337_ ) );
DFF_X1 \IFU/_602_ ( .D(\IFU/_379_ ), .CK(clock ), .Q(\_IFU_io_master_araddr [19] ), .QN(\IFU/_336_ ) );
DFF_X1 \IFU/_603_ ( .D(\IFU/_380_ ), .CK(clock ), .Q(\_IFU_io_master_araddr [20] ), .QN(\IFU/_335_ ) );
DFF_X1 \IFU/_604_ ( .D(\IFU/_381_ ), .CK(clock ), .Q(\_IFU_io_master_araddr [21] ), .QN(\IFU/_334_ ) );
DFF_X1 \IFU/_605_ ( .D(\IFU/_382_ ), .CK(clock ), .Q(\_IFU_io_master_araddr [22] ), .QN(\IFU/_333_ ) );
DFF_X1 \IFU/_606_ ( .D(\IFU/_383_ ), .CK(clock ), .Q(\_IFU_io_master_araddr [23] ), .QN(\IFU/_332_ ) );
DFF_X1 \IFU/_607_ ( .D(\IFU/_384_ ), .CK(clock ), .Q(\_IFU_io_master_araddr [24] ), .QN(\IFU/_331_ ) );
DFF_X1 \IFU/_608_ ( .D(\IFU/_385_ ), .CK(clock ), .Q(\_IFU_io_master_araddr [25] ), .QN(\IFU/_330_ ) );
DFF_X1 \IFU/_609_ ( .D(\IFU/_386_ ), .CK(clock ), .Q(\_IFU_io_master_araddr [26] ), .QN(\IFU/_329_ ) );
DFF_X1 \IFU/_610_ ( .D(\IFU/_387_ ), .CK(clock ), .Q(\_IFU_io_master_araddr [27] ), .QN(\IFU/_328_ ) );
DFF_X1 \IFU/_611_ ( .D(\IFU/_388_ ), .CK(clock ), .Q(\_IFU_io_master_araddr [28] ), .QN(\IFU/_327_ ) );
DFF_X1 \IFU/_612_ ( .D(\IFU/_389_ ), .CK(clock ), .Q(\_IFU_io_master_araddr [29] ), .QN(\IFU/_326_ ) );
DFF_X1 \IFU/_613_ ( .D(\IFU/_390_ ), .CK(clock ), .Q(\_IFU_io_master_araddr [30] ), .QN(\IFU/_325_ ) );
DFF_X1 \IFU/_614_ ( .D(\IFU/_391_ ), .CK(clock ), .Q(\_IFU_io_master_araddr [31] ), .QN(\IFU/_324_ ) );
DFF_X1 \IFU/_615_ ( .D(\IFU/_392_ ), .CK(clock ), .Q(\_IFU_io_out_bits_instruction [0] ), .QN(\IFU/_323_ ) );
DFF_X1 \IFU/_616_ ( .D(\IFU/_393_ ), .CK(clock ), .Q(\_IFU_io_out_bits_instruction [1] ), .QN(\IFU/_322_ ) );
DFF_X1 \IFU/_617_ ( .D(\IFU/_394_ ), .CK(clock ), .Q(\_IFU_io_out_bits_instruction [2] ), .QN(\IFU/_321_ ) );
DFF_X1 \IFU/_618_ ( .D(\IFU/_395_ ), .CK(clock ), .Q(\_IFU_io_out_bits_instruction [3] ), .QN(\IFU/_320_ ) );
DFF_X1 \IFU/_619_ ( .D(\IFU/_396_ ), .CK(clock ), .Q(\_IFU_io_out_bits_instruction [4] ), .QN(\IFU/_319_ ) );
DFF_X1 \IFU/_620_ ( .D(\IFU/_397_ ), .CK(clock ), .Q(\_IFU_io_out_bits_instruction [5] ), .QN(\IFU/_318_ ) );
DFF_X1 \IFU/_621_ ( .D(\IFU/_398_ ), .CK(clock ), .Q(\_IFU_io_out_bits_instruction [6] ), .QN(\IFU/_317_ ) );
DFF_X1 \IFU/_622_ ( .D(\IFU/_399_ ), .CK(clock ), .Q(\_IFU_io_out_bits_instruction [7] ), .QN(\IFU/_316_ ) );
DFF_X1 \IFU/_623_ ( .D(\IFU/_400_ ), .CK(clock ), .Q(\_IFU_io_out_bits_instruction [8] ), .QN(\IFU/_315_ ) );
DFF_X1 \IFU/_624_ ( .D(\IFU/_401_ ), .CK(clock ), .Q(\_IFU_io_out_bits_instruction [9] ), .QN(\IFU/_314_ ) );
DFF_X1 \IFU/_625_ ( .D(\IFU/_402_ ), .CK(clock ), .Q(\_IFU_io_out_bits_instruction [10] ), .QN(\IFU/_313_ ) );
DFF_X1 \IFU/_626_ ( .D(\IFU/_403_ ), .CK(clock ), .Q(\_IFU_io_out_bits_instruction [11] ), .QN(\IFU/_312_ ) );
DFF_X1 \IFU/_627_ ( .D(\IFU/_404_ ), .CK(clock ), .Q(\_IFU_io_out_bits_instruction [12] ), .QN(\IFU/_311_ ) );
DFF_X1 \IFU/_628_ ( .D(\IFU/_405_ ), .CK(clock ), .Q(\_IFU_io_out_bits_instruction [13] ), .QN(\IFU/_310_ ) );
DFF_X1 \IFU/_629_ ( .D(\IFU/_406_ ), .CK(clock ), .Q(\_IFU_io_out_bits_instruction [14] ), .QN(\IFU/_309_ ) );
DFF_X1 \IFU/_630_ ( .D(\IFU/_407_ ), .CK(clock ), .Q(\_IFU_io_out_bits_instruction [15] ), .QN(\IFU/_308_ ) );
DFF_X1 \IFU/_631_ ( .D(\IFU/_408_ ), .CK(clock ), .Q(\_IFU_io_out_bits_instruction [16] ), .QN(\IFU/_307_ ) );
DFF_X1 \IFU/_632_ ( .D(\IFU/_409_ ), .CK(clock ), .Q(\_IFU_io_out_bits_instruction [17] ), .QN(\IFU/_306_ ) );
DFF_X1 \IFU/_633_ ( .D(\IFU/_410_ ), .CK(clock ), .Q(\_IFU_io_out_bits_instruction [18] ), .QN(\IFU/_305_ ) );
DFF_X1 \IFU/_634_ ( .D(\IFU/_411_ ), .CK(clock ), .Q(\_IFU_io_out_bits_instruction [19] ), .QN(\IFU/_304_ ) );
DFF_X1 \IFU/_635_ ( .D(\IFU/_412_ ), .CK(clock ), .Q(\_IFU_io_out_bits_instruction [20] ), .QN(\IFU/_303_ ) );
DFF_X1 \IFU/_636_ ( .D(\IFU/_413_ ), .CK(clock ), .Q(\_IFU_io_out_bits_instruction [21] ), .QN(\IFU/_302_ ) );
DFF_X1 \IFU/_637_ ( .D(\IFU/_414_ ), .CK(clock ), .Q(\_IFU_io_out_bits_instruction [22] ), .QN(\IFU/_301_ ) );
DFF_X1 \IFU/_638_ ( .D(\IFU/_415_ ), .CK(clock ), .Q(\_IFU_io_out_bits_instruction [23] ), .QN(\IFU/_300_ ) );
DFF_X1 \IFU/_639_ ( .D(\IFU/_416_ ), .CK(clock ), .Q(\_IFU_io_out_bits_instruction [24] ), .QN(\IFU/_299_ ) );
DFF_X1 \IFU/_640_ ( .D(\IFU/_417_ ), .CK(clock ), .Q(\_IFU_io_out_bits_instruction [25] ), .QN(\IFU/_298_ ) );
DFF_X1 \IFU/_641_ ( .D(\IFU/_418_ ), .CK(clock ), .Q(\_IFU_io_out_bits_instruction [26] ), .QN(\IFU/_297_ ) );
DFF_X1 \IFU/_642_ ( .D(\IFU/_419_ ), .CK(clock ), .Q(\_IFU_io_out_bits_instruction [27] ), .QN(\IFU/_296_ ) );
DFF_X1 \IFU/_643_ ( .D(\IFU/_420_ ), .CK(clock ), .Q(\_IFU_io_out_bits_instruction [28] ), .QN(\IFU/_295_ ) );
DFF_X1 \IFU/_644_ ( .D(\IFU/_421_ ), .CK(clock ), .Q(\_IFU_io_out_bits_instruction [29] ), .QN(\IFU/_294_ ) );
DFF_X1 \IFU/_645_ ( .D(\IFU/_422_ ), .CK(clock ), .Q(\_IFU_io_out_bits_instruction [30] ), .QN(\IFU/_293_ ) );
DFF_X1 \IFU/_646_ ( .D(\IFU/_423_ ), .CK(clock ), .Q(\_IFU_io_out_bits_instruction [31] ), .QN(\IFU/_292_ ) );
BUF_X1 \IFU/_647_ ( .A(\_IFU_io_master_araddr [0] ), .Z(\_IFU_io_out_bits_pc [0] ) );
BUF_X1 \IFU/_648_ ( .A(\_IFU_io_master_araddr [1] ), .Z(\_IFU_io_out_bits_pc [1] ) );
BUF_X1 \IFU/_649_ ( .A(\_IFU_io_master_araddr [2] ), .Z(\_IFU_io_out_bits_pc [2] ) );
BUF_X1 \IFU/_650_ ( .A(\_IFU_io_master_araddr [3] ), .Z(\_IFU_io_out_bits_pc [3] ) );
BUF_X1 \IFU/_651_ ( .A(\_IFU_io_master_araddr [4] ), .Z(\_IFU_io_out_bits_pc [4] ) );
BUF_X1 \IFU/_652_ ( .A(\_IFU_io_master_araddr [5] ), .Z(\_IFU_io_out_bits_pc [5] ) );
BUF_X1 \IFU/_653_ ( .A(\_IFU_io_master_araddr [6] ), .Z(\_IFU_io_out_bits_pc [6] ) );
BUF_X1 \IFU/_654_ ( .A(\_IFU_io_master_araddr [7] ), .Z(\_IFU_io_out_bits_pc [7] ) );
BUF_X1 \IFU/_655_ ( .A(\_IFU_io_master_araddr [8] ), .Z(\_IFU_io_out_bits_pc [8] ) );
BUF_X1 \IFU/_656_ ( .A(\_IFU_io_master_araddr [9] ), .Z(\_IFU_io_out_bits_pc [9] ) );
BUF_X1 \IFU/_657_ ( .A(\_IFU_io_master_araddr [10] ), .Z(\_IFU_io_out_bits_pc [10] ) );
BUF_X1 \IFU/_658_ ( .A(\_IFU_io_master_araddr [11] ), .Z(\_IFU_io_out_bits_pc [11] ) );
BUF_X1 \IFU/_659_ ( .A(\_IFU_io_master_araddr [12] ), .Z(\_IFU_io_out_bits_pc [12] ) );
BUF_X1 \IFU/_660_ ( .A(\_IFU_io_master_araddr [13] ), .Z(\_IFU_io_out_bits_pc [13] ) );
BUF_X1 \IFU/_661_ ( .A(\_IFU_io_master_araddr [14] ), .Z(\_IFU_io_out_bits_pc [14] ) );
BUF_X1 \IFU/_662_ ( .A(\_IFU_io_master_araddr [15] ), .Z(\_IFU_io_out_bits_pc [15] ) );
BUF_X1 \IFU/_663_ ( .A(\_IFU_io_master_araddr [16] ), .Z(\_IFU_io_out_bits_pc [16] ) );
BUF_X1 \IFU/_664_ ( .A(\_IFU_io_master_araddr [17] ), .Z(\_IFU_io_out_bits_pc [17] ) );
BUF_X1 \IFU/_665_ ( .A(\_IFU_io_master_araddr [18] ), .Z(\_IFU_io_out_bits_pc [18] ) );
BUF_X1 \IFU/_666_ ( .A(\_IFU_io_master_araddr [19] ), .Z(\_IFU_io_out_bits_pc [19] ) );
BUF_X1 \IFU/_667_ ( .A(\_IFU_io_master_araddr [20] ), .Z(\_IFU_io_out_bits_pc [20] ) );
BUF_X1 \IFU/_668_ ( .A(\_IFU_io_master_araddr [21] ), .Z(\_IFU_io_out_bits_pc [21] ) );
BUF_X1 \IFU/_669_ ( .A(\_IFU_io_master_araddr [22] ), .Z(\_IFU_io_out_bits_pc [22] ) );
BUF_X1 \IFU/_670_ ( .A(\_IFU_io_master_araddr [23] ), .Z(\_IFU_io_out_bits_pc [23] ) );
BUF_X1 \IFU/_671_ ( .A(\_IFU_io_master_araddr [24] ), .Z(\_IFU_io_out_bits_pc [24] ) );
BUF_X1 \IFU/_672_ ( .A(\_IFU_io_master_araddr [25] ), .Z(\_IFU_io_out_bits_pc [25] ) );
BUF_X1 \IFU/_673_ ( .A(\_IFU_io_master_araddr [26] ), .Z(\_IFU_io_out_bits_pc [26] ) );
BUF_X1 \IFU/_674_ ( .A(\_IFU_io_master_araddr [27] ), .Z(\_IFU_io_out_bits_pc [27] ) );
BUF_X1 \IFU/_675_ ( .A(\_IFU_io_master_araddr [28] ), .Z(\_IFU_io_out_bits_pc [28] ) );
BUF_X1 \IFU/_676_ ( .A(\_IFU_io_master_araddr [29] ), .Z(\_IFU_io_out_bits_pc [29] ) );
BUF_X1 \IFU/_677_ ( .A(\_IFU_io_master_araddr [30] ), .Z(\_IFU_io_out_bits_pc [30] ) );
BUF_X1 \IFU/_678_ ( .A(\_IFU_io_master_araddr [31] ), .Z(\_IFU_io_out_bits_pc [31] ) );
BUF_X1 \IFU/_679_ ( .A(\IFU/state [0] ), .Z(\IFU/_290_ ) );
BUF_X1 \IFU/_680_ ( .A(\IFU/state [1] ), .Z(\IFU/_291_ ) );
BUF_X1 \IFU/_681_ ( .A(\IFU/_201_ ), .Z(_IFU_io_out_valid ) );
BUF_X1 \IFU/_682_ ( .A(\IFU/_166_ ), .Z(_IFU_io_master_rready ) );
BUF_X1 \IFU/_683_ ( .A(\IFU/_133_ ), .Z(_IFU_io_master_arvalid ) );
BUF_X1 \IFU/_684_ ( .A(\IFU/_098_ ), .Z(_IFU_io_in_ready ) );
BUF_X1 \IFU/_685_ ( .A(_IDU_io_in_ready ), .Z(\IFU/_200_ ) );
BUF_X1 \IFU/_686_ ( .A(_AXI4Interconnect_io_fanIn_0_rvalid ), .Z(\IFU/_167_ ) );
BUF_X1 \IFU/_687_ ( .A(_AXI4Interconnect_io_fanIn_0_arready ), .Z(\IFU/_132_ ) );
BUF_X1 \IFU/_688_ ( .A(_WBU_io_out_valid ), .Z(\IFU/_099_ ) );
BUF_X1 \IFU/_689_ ( .A(\_IFU_io_master_araddr [0] ), .Z(\IFU/_100_ ) );
BUF_X1 \IFU/_690_ ( .A(\_WBU_io_out_bits_nextPc [0] ), .Z(\IFU/_066_ ) );
BUF_X1 \IFU/_691_ ( .A(\_IFU_io_master_araddr [1] ), .Z(\IFU/_111_ ) );
BUF_X1 \IFU/_692_ ( .A(\_WBU_io_out_bits_nextPc [1] ), .Z(\IFU/_077_ ) );
BUF_X1 \IFU/_693_ ( .A(\_IFU_io_master_araddr [2] ), .Z(\IFU/_122_ ) );
BUF_X1 \IFU/_694_ ( .A(\_WBU_io_out_bits_nextPc [2] ), .Z(\IFU/_088_ ) );
BUF_X1 \IFU/_695_ ( .A(\_IFU_io_master_araddr [3] ), .Z(\IFU/_125_ ) );
BUF_X1 \IFU/_696_ ( .A(\_WBU_io_out_bits_nextPc [3] ), .Z(\IFU/_091_ ) );
BUF_X1 \IFU/_697_ ( .A(\_IFU_io_master_araddr [4] ), .Z(\IFU/_126_ ) );
BUF_X1 \IFU/_698_ ( .A(\_WBU_io_out_bits_nextPc [4] ), .Z(\IFU/_092_ ) );
BUF_X1 \IFU/_699_ ( .A(\_IFU_io_master_araddr [5] ), .Z(\IFU/_127_ ) );
BUF_X1 \IFU/_700_ ( .A(\_WBU_io_out_bits_nextPc [5] ), .Z(\IFU/_093_ ) );
BUF_X1 \IFU/_701_ ( .A(\_IFU_io_master_araddr [6] ), .Z(\IFU/_128_ ) );
BUF_X1 \IFU/_702_ ( .A(\_WBU_io_out_bits_nextPc [6] ), .Z(\IFU/_094_ ) );
BUF_X1 \IFU/_703_ ( .A(\_IFU_io_master_araddr [7] ), .Z(\IFU/_129_ ) );
BUF_X1 \IFU/_704_ ( .A(\_WBU_io_out_bits_nextPc [7] ), .Z(\IFU/_095_ ) );
BUF_X1 \IFU/_705_ ( .A(\_IFU_io_master_araddr [8] ), .Z(\IFU/_130_ ) );
BUF_X1 \IFU/_706_ ( .A(\_WBU_io_out_bits_nextPc [8] ), .Z(\IFU/_096_ ) );
BUF_X1 \IFU/_707_ ( .A(\_IFU_io_master_araddr [9] ), .Z(\IFU/_131_ ) );
BUF_X1 \IFU/_708_ ( .A(\_WBU_io_out_bits_nextPc [9] ), .Z(\IFU/_097_ ) );
BUF_X1 \IFU/_709_ ( .A(\_IFU_io_master_araddr [10] ), .Z(\IFU/_101_ ) );
BUF_X1 \IFU/_710_ ( .A(\_WBU_io_out_bits_nextPc [10] ), .Z(\IFU/_067_ ) );
BUF_X1 \IFU/_711_ ( .A(\_IFU_io_master_araddr [11] ), .Z(\IFU/_102_ ) );
BUF_X1 \IFU/_712_ ( .A(\_WBU_io_out_bits_nextPc [11] ), .Z(\IFU/_068_ ) );
BUF_X1 \IFU/_713_ ( .A(\_IFU_io_master_araddr [12] ), .Z(\IFU/_103_ ) );
BUF_X1 \IFU/_714_ ( .A(\_WBU_io_out_bits_nextPc [12] ), .Z(\IFU/_069_ ) );
BUF_X1 \IFU/_715_ ( .A(\_IFU_io_master_araddr [13] ), .Z(\IFU/_104_ ) );
BUF_X1 \IFU/_716_ ( .A(\_WBU_io_out_bits_nextPc [13] ), .Z(\IFU/_070_ ) );
BUF_X1 \IFU/_717_ ( .A(\_IFU_io_master_araddr [14] ), .Z(\IFU/_105_ ) );
BUF_X1 \IFU/_718_ ( .A(\_WBU_io_out_bits_nextPc [14] ), .Z(\IFU/_071_ ) );
BUF_X1 \IFU/_719_ ( .A(\_IFU_io_master_araddr [15] ), .Z(\IFU/_106_ ) );
BUF_X1 \IFU/_720_ ( .A(\_WBU_io_out_bits_nextPc [15] ), .Z(\IFU/_072_ ) );
BUF_X1 \IFU/_721_ ( .A(\_IFU_io_master_araddr [16] ), .Z(\IFU/_107_ ) );
BUF_X1 \IFU/_722_ ( .A(\_WBU_io_out_bits_nextPc [16] ), .Z(\IFU/_073_ ) );
BUF_X1 \IFU/_723_ ( .A(\_IFU_io_master_araddr [17] ), .Z(\IFU/_108_ ) );
BUF_X1 \IFU/_724_ ( .A(\_WBU_io_out_bits_nextPc [17] ), .Z(\IFU/_074_ ) );
BUF_X1 \IFU/_725_ ( .A(\_IFU_io_master_araddr [18] ), .Z(\IFU/_109_ ) );
BUF_X1 \IFU/_726_ ( .A(\_WBU_io_out_bits_nextPc [18] ), .Z(\IFU/_075_ ) );
BUF_X1 \IFU/_727_ ( .A(\_IFU_io_master_araddr [19] ), .Z(\IFU/_110_ ) );
BUF_X1 \IFU/_728_ ( .A(\_WBU_io_out_bits_nextPc [19] ), .Z(\IFU/_076_ ) );
BUF_X1 \IFU/_729_ ( .A(\_IFU_io_master_araddr [20] ), .Z(\IFU/_112_ ) );
BUF_X1 \IFU/_730_ ( .A(\_WBU_io_out_bits_nextPc [20] ), .Z(\IFU/_078_ ) );
BUF_X1 \IFU/_731_ ( .A(\_IFU_io_master_araddr [21] ), .Z(\IFU/_113_ ) );
BUF_X1 \IFU/_732_ ( .A(\_WBU_io_out_bits_nextPc [21] ), .Z(\IFU/_079_ ) );
BUF_X1 \IFU/_733_ ( .A(\_IFU_io_master_araddr [22] ), .Z(\IFU/_114_ ) );
BUF_X1 \IFU/_734_ ( .A(\_WBU_io_out_bits_nextPc [22] ), .Z(\IFU/_080_ ) );
BUF_X1 \IFU/_735_ ( .A(\_IFU_io_master_araddr [23] ), .Z(\IFU/_115_ ) );
BUF_X1 \IFU/_736_ ( .A(\_WBU_io_out_bits_nextPc [23] ), .Z(\IFU/_081_ ) );
BUF_X1 \IFU/_737_ ( .A(\_IFU_io_master_araddr [24] ), .Z(\IFU/_116_ ) );
BUF_X1 \IFU/_738_ ( .A(\_WBU_io_out_bits_nextPc [24] ), .Z(\IFU/_082_ ) );
BUF_X1 \IFU/_739_ ( .A(\_IFU_io_master_araddr [25] ), .Z(\IFU/_117_ ) );
BUF_X1 \IFU/_740_ ( .A(\_WBU_io_out_bits_nextPc [25] ), .Z(\IFU/_083_ ) );
BUF_X1 \IFU/_741_ ( .A(\_IFU_io_master_araddr [26] ), .Z(\IFU/_118_ ) );
BUF_X1 \IFU/_742_ ( .A(\_WBU_io_out_bits_nextPc [26] ), .Z(\IFU/_084_ ) );
BUF_X1 \IFU/_743_ ( .A(\_IFU_io_master_araddr [27] ), .Z(\IFU/_119_ ) );
BUF_X1 \IFU/_744_ ( .A(\_WBU_io_out_bits_nextPc [27] ), .Z(\IFU/_085_ ) );
BUF_X1 \IFU/_745_ ( .A(\_IFU_io_master_araddr [28] ), .Z(\IFU/_120_ ) );
BUF_X1 \IFU/_746_ ( .A(\_WBU_io_out_bits_nextPc [28] ), .Z(\IFU/_086_ ) );
BUF_X1 \IFU/_747_ ( .A(\_IFU_io_master_araddr [29] ), .Z(\IFU/_121_ ) );
BUF_X1 \IFU/_748_ ( .A(\_WBU_io_out_bits_nextPc [29] ), .Z(\IFU/_087_ ) );
BUF_X1 \IFU/_749_ ( .A(\_IFU_io_master_araddr [30] ), .Z(\IFU/_123_ ) );
BUF_X1 \IFU/_750_ ( .A(\_WBU_io_out_bits_nextPc [30] ), .Z(\IFU/_089_ ) );
BUF_X1 \IFU/_751_ ( .A(\_IFU_io_master_araddr [31] ), .Z(\IFU/_124_ ) );
BUF_X1 \IFU/_752_ ( .A(\_WBU_io_out_bits_nextPc [31] ), .Z(\IFU/_090_ ) );
BUF_X1 \IFU/_753_ ( .A(\_IFU_io_out_bits_instruction [0] ), .Z(\IFU/_168_ ) );
BUF_X1 \IFU/_754_ ( .A(\_AXI4Interconnect_io_fanIn_0_rdata [0] ), .Z(\IFU/_134_ ) );
BUF_X1 \IFU/_755_ ( .A(\_IFU_io_out_bits_instruction [1] ), .Z(\IFU/_179_ ) );
BUF_X1 \IFU/_756_ ( .A(\_AXI4Interconnect_io_fanIn_0_rdata [1] ), .Z(\IFU/_145_ ) );
BUF_X1 \IFU/_757_ ( .A(\_IFU_io_out_bits_instruction [2] ), .Z(\IFU/_190_ ) );
BUF_X1 \IFU/_758_ ( .A(\_AXI4Interconnect_io_fanIn_0_rdata [2] ), .Z(\IFU/_156_ ) );
BUF_X1 \IFU/_759_ ( .A(\_IFU_io_out_bits_instruction [3] ), .Z(\IFU/_193_ ) );
BUF_X1 \IFU/_760_ ( .A(\_AXI4Interconnect_io_fanIn_0_rdata [3] ), .Z(\IFU/_159_ ) );
BUF_X1 \IFU/_761_ ( .A(\_IFU_io_out_bits_instruction [4] ), .Z(\IFU/_194_ ) );
BUF_X1 \IFU/_762_ ( .A(\_AXI4Interconnect_io_fanIn_0_rdata [4] ), .Z(\IFU/_160_ ) );
BUF_X1 \IFU/_763_ ( .A(\_IFU_io_out_bits_instruction [5] ), .Z(\IFU/_195_ ) );
BUF_X1 \IFU/_764_ ( .A(\_AXI4Interconnect_io_fanIn_0_rdata [5] ), .Z(\IFU/_161_ ) );
BUF_X1 \IFU/_765_ ( .A(\_IFU_io_out_bits_instruction [6] ), .Z(\IFU/_196_ ) );
BUF_X1 \IFU/_766_ ( .A(\_AXI4Interconnect_io_fanIn_0_rdata [6] ), .Z(\IFU/_162_ ) );
BUF_X1 \IFU/_767_ ( .A(\_IFU_io_out_bits_instruction [7] ), .Z(\IFU/_197_ ) );
BUF_X1 \IFU/_768_ ( .A(\_AXI4Interconnect_io_fanIn_0_rdata [7] ), .Z(\IFU/_163_ ) );
BUF_X1 \IFU/_769_ ( .A(\_IFU_io_out_bits_instruction [8] ), .Z(\IFU/_198_ ) );
BUF_X1 \IFU/_770_ ( .A(\_AXI4Interconnect_io_fanIn_0_rdata [8] ), .Z(\IFU/_164_ ) );
BUF_X1 \IFU/_771_ ( .A(\_IFU_io_out_bits_instruction [9] ), .Z(\IFU/_199_ ) );
BUF_X1 \IFU/_772_ ( .A(\_AXI4Interconnect_io_fanIn_0_rdata [9] ), .Z(\IFU/_165_ ) );
BUF_X1 \IFU/_773_ ( .A(\_IFU_io_out_bits_instruction [10] ), .Z(\IFU/_169_ ) );
BUF_X1 \IFU/_774_ ( .A(\_AXI4Interconnect_io_fanIn_0_rdata [10] ), .Z(\IFU/_135_ ) );
BUF_X1 \IFU/_775_ ( .A(\_IFU_io_out_bits_instruction [11] ), .Z(\IFU/_170_ ) );
BUF_X1 \IFU/_776_ ( .A(\_AXI4Interconnect_io_fanIn_0_rdata [11] ), .Z(\IFU/_136_ ) );
BUF_X1 \IFU/_777_ ( .A(\_IFU_io_out_bits_instruction [12] ), .Z(\IFU/_171_ ) );
BUF_X1 \IFU/_778_ ( .A(\_AXI4Interconnect_io_fanIn_0_rdata [12] ), .Z(\IFU/_137_ ) );
BUF_X1 \IFU/_779_ ( .A(\_IFU_io_out_bits_instruction [13] ), .Z(\IFU/_172_ ) );
BUF_X1 \IFU/_780_ ( .A(\_AXI4Interconnect_io_fanIn_0_rdata [13] ), .Z(\IFU/_138_ ) );
BUF_X1 \IFU/_781_ ( .A(\_IFU_io_out_bits_instruction [14] ), .Z(\IFU/_173_ ) );
BUF_X1 \IFU/_782_ ( .A(\_AXI4Interconnect_io_fanIn_0_rdata [14] ), .Z(\IFU/_139_ ) );
BUF_X1 \IFU/_783_ ( .A(\_IFU_io_out_bits_instruction [15] ), .Z(\IFU/_174_ ) );
BUF_X1 \IFU/_784_ ( .A(\_AXI4Interconnect_io_fanIn_0_rdata [15] ), .Z(\IFU/_140_ ) );
BUF_X1 \IFU/_785_ ( .A(\_IFU_io_out_bits_instruction [16] ), .Z(\IFU/_175_ ) );
BUF_X1 \IFU/_786_ ( .A(\_AXI4Interconnect_io_fanIn_0_rdata [16] ), .Z(\IFU/_141_ ) );
BUF_X1 \IFU/_787_ ( .A(\_IFU_io_out_bits_instruction [17] ), .Z(\IFU/_176_ ) );
BUF_X1 \IFU/_788_ ( .A(\_AXI4Interconnect_io_fanIn_0_rdata [17] ), .Z(\IFU/_142_ ) );
BUF_X1 \IFU/_789_ ( .A(\_IFU_io_out_bits_instruction [18] ), .Z(\IFU/_177_ ) );
BUF_X1 \IFU/_790_ ( .A(\_AXI4Interconnect_io_fanIn_0_rdata [18] ), .Z(\IFU/_143_ ) );
BUF_X1 \IFU/_791_ ( .A(\_IFU_io_out_bits_instruction [19] ), .Z(\IFU/_178_ ) );
BUF_X1 \IFU/_792_ ( .A(\_AXI4Interconnect_io_fanIn_0_rdata [19] ), .Z(\IFU/_144_ ) );
BUF_X1 \IFU/_793_ ( .A(\_IFU_io_out_bits_instruction [20] ), .Z(\IFU/_180_ ) );
BUF_X1 \IFU/_794_ ( .A(\_AXI4Interconnect_io_fanIn_0_rdata [20] ), .Z(\IFU/_146_ ) );
BUF_X1 \IFU/_795_ ( .A(\_IFU_io_out_bits_instruction [21] ), .Z(\IFU/_181_ ) );
BUF_X1 \IFU/_796_ ( .A(\_AXI4Interconnect_io_fanIn_0_rdata [21] ), .Z(\IFU/_147_ ) );
BUF_X1 \IFU/_797_ ( .A(\_IFU_io_out_bits_instruction [22] ), .Z(\IFU/_182_ ) );
BUF_X1 \IFU/_798_ ( .A(\_AXI4Interconnect_io_fanIn_0_rdata [22] ), .Z(\IFU/_148_ ) );
BUF_X1 \IFU/_799_ ( .A(\_IFU_io_out_bits_instruction [23] ), .Z(\IFU/_183_ ) );
BUF_X1 \IFU/_800_ ( .A(\_AXI4Interconnect_io_fanIn_0_rdata [23] ), .Z(\IFU/_149_ ) );
BUF_X1 \IFU/_801_ ( .A(\_IFU_io_out_bits_instruction [24] ), .Z(\IFU/_184_ ) );
BUF_X1 \IFU/_802_ ( .A(\_AXI4Interconnect_io_fanIn_0_rdata [24] ), .Z(\IFU/_150_ ) );
BUF_X1 \IFU/_803_ ( .A(\_IFU_io_out_bits_instruction [25] ), .Z(\IFU/_185_ ) );
BUF_X1 \IFU/_804_ ( .A(\_AXI4Interconnect_io_fanIn_0_rdata [25] ), .Z(\IFU/_151_ ) );
BUF_X1 \IFU/_805_ ( .A(\_IFU_io_out_bits_instruction [26] ), .Z(\IFU/_186_ ) );
BUF_X1 \IFU/_806_ ( .A(\_AXI4Interconnect_io_fanIn_0_rdata [26] ), .Z(\IFU/_152_ ) );
BUF_X1 \IFU/_807_ ( .A(\_IFU_io_out_bits_instruction [27] ), .Z(\IFU/_187_ ) );
BUF_X1 \IFU/_808_ ( .A(\_AXI4Interconnect_io_fanIn_0_rdata [27] ), .Z(\IFU/_153_ ) );
BUF_X1 \IFU/_809_ ( .A(\_IFU_io_out_bits_instruction [28] ), .Z(\IFU/_188_ ) );
BUF_X1 \IFU/_810_ ( .A(\_AXI4Interconnect_io_fanIn_0_rdata [28] ), .Z(\IFU/_154_ ) );
BUF_X1 \IFU/_811_ ( .A(\_IFU_io_out_bits_instruction [29] ), .Z(\IFU/_189_ ) );
BUF_X1 \IFU/_812_ ( .A(\_AXI4Interconnect_io_fanIn_0_rdata [29] ), .Z(\IFU/_155_ ) );
BUF_X1 \IFU/_813_ ( .A(\_IFU_io_out_bits_instruction [30] ), .Z(\IFU/_191_ ) );
BUF_X1 \IFU/_814_ ( .A(\_AXI4Interconnect_io_fanIn_0_rdata [30] ), .Z(\IFU/_157_ ) );
BUF_X1 \IFU/_815_ ( .A(\_IFU_io_out_bits_instruction [31] ), .Z(\IFU/_192_ ) );
BUF_X1 \IFU/_816_ ( .A(\_AXI4Interconnect_io_fanIn_0_rdata [31] ), .Z(\IFU/_158_ ) );
BUF_X1 \IFU/_817_ ( .A(reset ), .Z(\IFU/_289_ ) );
BUF_X1 \IFU/_818_ ( .A(\IFU/_000_ ), .Z(\IFU/_358_ ) );
BUF_X1 \IFU/_819_ ( .A(\IFU/_001_ ), .Z(\IFU/_359_ ) );
BUF_X1 \IFU/_820_ ( .A(\IFU/_002_ ), .Z(\IFU/_360_ ) );
BUF_X1 \IFU/_821_ ( .A(\IFU/_003_ ), .Z(\IFU/_361_ ) );
BUF_X1 \IFU/_822_ ( .A(\IFU/_004_ ), .Z(\IFU/_362_ ) );
BUF_X1 \IFU/_823_ ( .A(\IFU/_005_ ), .Z(\IFU/_363_ ) );
BUF_X1 \IFU/_824_ ( .A(\IFU/_006_ ), .Z(\IFU/_364_ ) );
BUF_X1 \IFU/_825_ ( .A(\IFU/_007_ ), .Z(\IFU/_365_ ) );
BUF_X1 \IFU/_826_ ( .A(\IFU/_008_ ), .Z(\IFU/_366_ ) );
BUF_X1 \IFU/_827_ ( .A(\IFU/_009_ ), .Z(\IFU/_367_ ) );
BUF_X1 \IFU/_828_ ( .A(\IFU/_010_ ), .Z(\IFU/_368_ ) );
BUF_X1 \IFU/_829_ ( .A(\IFU/_011_ ), .Z(\IFU/_369_ ) );
BUF_X1 \IFU/_830_ ( .A(\IFU/_012_ ), .Z(\IFU/_370_ ) );
BUF_X1 \IFU/_831_ ( .A(\IFU/_013_ ), .Z(\IFU/_371_ ) );
BUF_X1 \IFU/_832_ ( .A(\IFU/_014_ ), .Z(\IFU/_372_ ) );
BUF_X1 \IFU/_833_ ( .A(\IFU/_015_ ), .Z(\IFU/_373_ ) );
BUF_X1 \IFU/_834_ ( .A(\IFU/_016_ ), .Z(\IFU/_374_ ) );
BUF_X1 \IFU/_835_ ( .A(\IFU/_017_ ), .Z(\IFU/_375_ ) );
BUF_X1 \IFU/_836_ ( .A(\IFU/_018_ ), .Z(\IFU/_376_ ) );
BUF_X1 \IFU/_837_ ( .A(\IFU/_019_ ), .Z(\IFU/_377_ ) );
BUF_X1 \IFU/_838_ ( .A(\IFU/_020_ ), .Z(\IFU/_378_ ) );
BUF_X1 \IFU/_839_ ( .A(\IFU/_021_ ), .Z(\IFU/_379_ ) );
BUF_X1 \IFU/_840_ ( .A(\IFU/_022_ ), .Z(\IFU/_380_ ) );
BUF_X1 \IFU/_841_ ( .A(\IFU/_023_ ), .Z(\IFU/_381_ ) );
BUF_X1 \IFU/_842_ ( .A(\IFU/_024_ ), .Z(\IFU/_382_ ) );
BUF_X1 \IFU/_843_ ( .A(\IFU/_025_ ), .Z(\IFU/_383_ ) );
BUF_X1 \IFU/_844_ ( .A(\IFU/_026_ ), .Z(\IFU/_384_ ) );
BUF_X1 \IFU/_845_ ( .A(\IFU/_027_ ), .Z(\IFU/_385_ ) );
BUF_X1 \IFU/_846_ ( .A(\IFU/_028_ ), .Z(\IFU/_386_ ) );
BUF_X1 \IFU/_847_ ( .A(\IFU/_029_ ), .Z(\IFU/_387_ ) );
BUF_X1 \IFU/_848_ ( .A(\IFU/_030_ ), .Z(\IFU/_388_ ) );
BUF_X1 \IFU/_849_ ( .A(\IFU/_031_ ), .Z(\IFU/_389_ ) );
BUF_X1 \IFU/_850_ ( .A(\IFU/_032_ ), .Z(\IFU/_390_ ) );
BUF_X1 \IFU/_851_ ( .A(\IFU/_033_ ), .Z(\IFU/_391_ ) );
BUF_X1 \IFU/_852_ ( .A(\IFU/_034_ ), .Z(\IFU/_392_ ) );
BUF_X1 \IFU/_853_ ( .A(\IFU/_035_ ), .Z(\IFU/_393_ ) );
BUF_X1 \IFU/_854_ ( .A(\IFU/_036_ ), .Z(\IFU/_394_ ) );
BUF_X1 \IFU/_855_ ( .A(\IFU/_037_ ), .Z(\IFU/_395_ ) );
BUF_X1 \IFU/_856_ ( .A(\IFU/_038_ ), .Z(\IFU/_396_ ) );
BUF_X1 \IFU/_857_ ( .A(\IFU/_039_ ), .Z(\IFU/_397_ ) );
BUF_X1 \IFU/_858_ ( .A(\IFU/_040_ ), .Z(\IFU/_398_ ) );
BUF_X1 \IFU/_859_ ( .A(\IFU/_041_ ), .Z(\IFU/_399_ ) );
BUF_X1 \IFU/_860_ ( .A(\IFU/_042_ ), .Z(\IFU/_400_ ) );
BUF_X1 \IFU/_861_ ( .A(\IFU/_043_ ), .Z(\IFU/_401_ ) );
BUF_X1 \IFU/_862_ ( .A(\IFU/_044_ ), .Z(\IFU/_402_ ) );
BUF_X1 \IFU/_863_ ( .A(\IFU/_045_ ), .Z(\IFU/_403_ ) );
BUF_X1 \IFU/_864_ ( .A(\IFU/_046_ ), .Z(\IFU/_404_ ) );
BUF_X1 \IFU/_865_ ( .A(\IFU/_047_ ), .Z(\IFU/_405_ ) );
BUF_X1 \IFU/_866_ ( .A(\IFU/_048_ ), .Z(\IFU/_406_ ) );
BUF_X1 \IFU/_867_ ( .A(\IFU/_049_ ), .Z(\IFU/_407_ ) );
BUF_X1 \IFU/_868_ ( .A(\IFU/_050_ ), .Z(\IFU/_408_ ) );
BUF_X1 \IFU/_869_ ( .A(\IFU/_051_ ), .Z(\IFU/_409_ ) );
BUF_X1 \IFU/_870_ ( .A(\IFU/_052_ ), .Z(\IFU/_410_ ) );
BUF_X1 \IFU/_871_ ( .A(\IFU/_053_ ), .Z(\IFU/_411_ ) );
BUF_X1 \IFU/_872_ ( .A(\IFU/_054_ ), .Z(\IFU/_412_ ) );
BUF_X1 \IFU/_873_ ( .A(\IFU/_055_ ), .Z(\IFU/_413_ ) );
BUF_X1 \IFU/_874_ ( .A(\IFU/_056_ ), .Z(\IFU/_414_ ) );
BUF_X1 \IFU/_875_ ( .A(\IFU/_057_ ), .Z(\IFU/_415_ ) );
BUF_X1 \IFU/_876_ ( .A(\IFU/_058_ ), .Z(\IFU/_416_ ) );
BUF_X1 \IFU/_877_ ( .A(\IFU/_059_ ), .Z(\IFU/_417_ ) );
BUF_X1 \IFU/_878_ ( .A(\IFU/_060_ ), .Z(\IFU/_418_ ) );
BUF_X1 \IFU/_879_ ( .A(\IFU/_061_ ), .Z(\IFU/_419_ ) );
BUF_X1 \IFU/_880_ ( .A(\IFU/_062_ ), .Z(\IFU/_420_ ) );
BUF_X1 \IFU/_881_ ( .A(\IFU/_063_ ), .Z(\IFU/_421_ ) );
BUF_X1 \IFU/_882_ ( .A(\IFU/_064_ ), .Z(\IFU/_422_ ) );
BUF_X1 \IFU/_883_ ( .A(\IFU/_065_ ), .Z(\IFU/_423_ ) );
INV_X1 \LSU/_0984_ ( .A(\LSU/_0005_ ), .ZN(\LSU/_0458_ ) );
AND3_X1 \LSU/_0985_ ( .A1(\LSU/_0458_ ), .A2(\LSU/_0718_ ), .A3(\LSU/_0717_ ), .ZN(\LSU/_0457_ ) );
INV_X32 \LSU/_0986_ ( .A(\LSU/_0718_ ), .ZN(\LSU/_0459_ ) );
AND3_X1 \LSU/_0987_ ( .A1(\LSU/_0459_ ), .A2(\LSU/_0717_ ), .A3(\LSU/_0719_ ), .ZN(\LSU/_0315_ ) );
NOR2_X4 \LSU/_0988_ ( .A1(\LSU/_0459_ ), .A2(\LSU/_0717_ ), .ZN(\LSU/_0460_ ) );
AND2_X2 \LSU/_0989_ ( .A1(\LSU/_0460_ ), .A2(\LSU/_0719_ ), .ZN(\LSU/_0384_ ) );
INV_X1 \LSU/_0990_ ( .A(\LSU/_0719_ ), .ZN(\LSU/_0461_ ) );
NOR3_X1 \LSU/_0991_ ( .A1(\LSU/_0461_ ), .A2(\LSU/_0718_ ), .A3(\LSU/_0717_ ), .ZN(\LSU/_0350_ ) );
NOR3_X1 \LSU/_0992_ ( .A1(\LSU/_0459_ ), .A2(\LSU/_0717_ ), .A3(\LSU/_0719_ ), .ZN(\LSU/_0462_ ) );
AND2_X1 \LSU/_0993_ ( .A1(\LSU/_0717_ ), .A2(\LSU/_0005_ ), .ZN(\LSU/_0463_ ) );
AOI21_X1 \LSU/_0994_ ( .A(\LSU/_0462_ ), .B1(\LSU/_0459_ ), .B2(\LSU/_0463_ ), .ZN(\LSU/_0464_ ) );
INV_X1 \LSU/_0995_ ( .A(\LSU/_0464_ ), .ZN(\LSU/_0349_ ) );
NOR3_X2 \LSU/_0996_ ( .A1(\LSU/_0458_ ), .A2(\LSU/_0718_ ), .A3(\LSU/_0717_ ), .ZN(\LSU/_0278_ ) );
INV_X1 \LSU/_0997_ ( .A(\LSU/_0717_ ), .ZN(\LSU/_0465_ ) );
NOR2_X1 \LSU/_0998_ ( .A1(\LSU/_0465_ ), .A2(\LSU/_0719_ ), .ZN(\LSU/_0418_ ) );
NOR2_X1 \LSU/_0999_ ( .A1(fanout_net_19 ), .A2(\LSU/_0327_ ), .ZN(\LSU/_0420_ ) );
INV_X32 \LSU/_1000_ ( .A(\LSU/_0314_ ), .ZN(\LSU/_0466_ ) );
INV_X32 \LSU/_1001_ ( .A(\LSU/_0313_ ), .ZN(\LSU/_0467_ ) );
NAND3_X1 \LSU/_1002_ ( .A1(\LSU/_0466_ ), .A2(\LSU/_0467_ ), .A3(\LSU/_0009_ ), .ZN(\LSU/_0468_ ) );
AND2_X1 \LSU/_1003_ ( .A1(\LSU/_0468_ ), .A2(\LSU/_0008_ ), .ZN(\LSU/_0421_ ) );
INV_X2 \LSU/_1004_ ( .A(fanout_net_19 ), .ZN(\LSU/_0469_ ) );
OAI21_X1 \LSU/_1005_ ( .A(\LSU/_0466_ ), .B1(\LSU/_0467_ ), .B2(\LSU/_0469_ ), .ZN(\LSU/_0470_ ) );
INV_X1 \LSU/_1006_ ( .A(\LSU/_0327_ ), .ZN(\LSU/_0471_ ) );
MUX2_X1 \LSU/_1007_ ( .A(\LSU/_0009_ ), .B(\LSU/_0470_ ), .S(\LSU/_0471_ ), .Z(\LSU/_0422_ ) );
NOR2_X4 \LSU/_1008_ ( .A1(\LSU/_0314_ ), .A2(\LSU/_0313_ ), .ZN(\LSU/_0472_ ) );
BUF_X4 \LSU/_1009_ ( .A(\LSU/_0472_ ), .Z(\LSU/_0473_ ) );
CLKBUF_X2 \LSU/_1010_ ( .A(\LSU/_0471_ ), .Z(\LSU/_0474_ ) );
AOI22_X1 \LSU/_1011_ ( .A1(\LSU/_0473_ ), .A2(\LSU/_0009_ ), .B1(\LSU/_0466_ ), .B2(\LSU/_0474_ ), .ZN(\LSU/_0423_ ) );
INV_X1 \LSU/_1012_ ( .A(\LSU/_0145_ ), .ZN(\LSU/_0475_ ) );
NOR3_X1 \LSU/_1013_ ( .A1(\LSU/_0475_ ), .A2(fanout_net_19 ), .A3(\LSU/_0327_ ), .ZN(\LSU/_0386_ ) );
INV_X1 \LSU/_1014_ ( .A(\LSU/_0156_ ), .ZN(\LSU/_0476_ ) );
NOR3_X1 \LSU/_1015_ ( .A1(\LSU/_0476_ ), .A2(fanout_net_19 ), .A3(\LSU/_0327_ ), .ZN(\LSU/_0397_ ) );
INV_X1 \LSU/_1016_ ( .A(\LSU/_0167_ ), .ZN(\LSU/_0477_ ) );
NOR3_X1 \LSU/_1017_ ( .A1(\LSU/_0477_ ), .A2(fanout_net_19 ), .A3(\LSU/_0327_ ), .ZN(\LSU/_0408_ ) );
INV_X1 \LSU/_1018_ ( .A(\LSU/_0170_ ), .ZN(\LSU/_0478_ ) );
NOR3_X1 \LSU/_1019_ ( .A1(\LSU/_0478_ ), .A2(fanout_net_19 ), .A3(\LSU/_0327_ ), .ZN(\LSU/_0411_ ) );
INV_X1 \LSU/_1020_ ( .A(\LSU/_0171_ ), .ZN(\LSU/_0479_ ) );
NOR3_X1 \LSU/_1021_ ( .A1(\LSU/_0479_ ), .A2(fanout_net_19 ), .A3(\LSU/_0327_ ), .ZN(\LSU/_0412_ ) );
INV_X1 \LSU/_1022_ ( .A(\LSU/_0172_ ), .ZN(\LSU/_0480_ ) );
NOR3_X1 \LSU/_1023_ ( .A1(\LSU/_0480_ ), .A2(fanout_net_19 ), .A3(\LSU/_0327_ ), .ZN(\LSU/_0413_ ) );
INV_X1 \LSU/_1024_ ( .A(\LSU/_0173_ ), .ZN(\LSU/_0481_ ) );
NOR3_X1 \LSU/_1025_ ( .A1(\LSU/_0481_ ), .A2(fanout_net_19 ), .A3(\LSU/_0327_ ), .ZN(\LSU/_0414_ ) );
INV_X1 \LSU/_1026_ ( .A(\LSU/_0174_ ), .ZN(\LSU/_0482_ ) );
NOR3_X1 \LSU/_1027_ ( .A1(\LSU/_0482_ ), .A2(fanout_net_19 ), .A3(\LSU/_0327_ ), .ZN(\LSU/_0415_ ) );
MUX2_X1 \LSU/_1028_ ( .A(\LSU/_0175_ ), .B(\LSU/_0145_ ), .S(fanout_net_19 ), .Z(\LSU/_0483_ ) );
AND2_X1 \LSU/_1029_ ( .A1(\LSU/_0483_ ), .A2(\LSU/_0474_ ), .ZN(\LSU/_0416_ ) );
MUX2_X1 \LSU/_1030_ ( .A(\LSU/_0176_ ), .B(\LSU/_0156_ ), .S(fanout_net_19 ), .Z(\LSU/_0484_ ) );
AND2_X1 \LSU/_1031_ ( .A1(\LSU/_0484_ ), .A2(\LSU/_0474_ ), .ZN(\LSU/_0417_ ) );
MUX2_X1 \LSU/_1032_ ( .A(\LSU/_0146_ ), .B(\LSU/_0167_ ), .S(fanout_net_19 ), .Z(\LSU/_0485_ ) );
AND2_X1 \LSU/_1033_ ( .A1(\LSU/_0485_ ), .A2(\LSU/_0474_ ), .ZN(\LSU/_0387_ ) );
MUX2_X1 \LSU/_1034_ ( .A(\LSU/_0147_ ), .B(\LSU/_0170_ ), .S(fanout_net_19 ), .Z(\LSU/_0486_ ) );
AND2_X1 \LSU/_1035_ ( .A1(\LSU/_0486_ ), .A2(\LSU/_0474_ ), .ZN(\LSU/_0388_ ) );
MUX2_X1 \LSU/_1036_ ( .A(\LSU/_0148_ ), .B(\LSU/_0171_ ), .S(fanout_net_19 ), .Z(\LSU/_0487_ ) );
AND2_X1 \LSU/_1037_ ( .A1(\LSU/_0487_ ), .A2(\LSU/_0474_ ), .ZN(\LSU/_0389_ ) );
MUX2_X1 \LSU/_1038_ ( .A(\LSU/_0149_ ), .B(\LSU/_0172_ ), .S(fanout_net_19 ), .Z(\LSU/_0488_ ) );
AND2_X1 \LSU/_1039_ ( .A1(\LSU/_0488_ ), .A2(\LSU/_0474_ ), .ZN(\LSU/_0390_ ) );
MUX2_X1 \LSU/_1040_ ( .A(\LSU/_0150_ ), .B(\LSU/_0173_ ), .S(fanout_net_19 ), .Z(\LSU/_0489_ ) );
AND2_X1 \LSU/_1041_ ( .A1(\LSU/_0489_ ), .A2(\LSU/_0474_ ), .ZN(\LSU/_0391_ ) );
MUX2_X1 \LSU/_1042_ ( .A(\LSU/_0151_ ), .B(\LSU/_0174_ ), .S(fanout_net_19 ), .Z(\LSU/_0490_ ) );
AND2_X1 \LSU/_1043_ ( .A1(\LSU/_0490_ ), .A2(\LSU/_0474_ ), .ZN(\LSU/_0392_ ) );
OAI21_X1 \LSU/_1044_ ( .A(\LSU/_0474_ ), .B1(\LSU/_0469_ ), .B2(\LSU/_0175_ ), .ZN(\LSU/_0491_ ) );
NOR2_X1 \LSU/_1045_ ( .A1(fanout_net_19 ), .A2(\LSU/_0152_ ), .ZN(\LSU/_0492_ ) );
NAND2_X1 \LSU/_1046_ ( .A1(\LSU/_0469_ ), .A2(\LSU/_0327_ ), .ZN(\LSU/_0493_ ) );
OAI22_X1 \LSU/_1047_ ( .A1(\LSU/_0491_ ), .A2(\LSU/_0492_ ), .B1(\LSU/_0493_ ), .B2(\LSU/_0475_ ), .ZN(\LSU/_0393_ ) );
OAI21_X1 \LSU/_1048_ ( .A(\LSU/_0471_ ), .B1(\LSU/_0469_ ), .B2(\LSU/_0176_ ), .ZN(\LSU/_0494_ ) );
NOR2_X1 \LSU/_1049_ ( .A1(fanout_net_19 ), .A2(\LSU/_0153_ ), .ZN(\LSU/_0495_ ) );
OAI22_X1 \LSU/_1050_ ( .A1(\LSU/_0494_ ), .A2(\LSU/_0495_ ), .B1(\LSU/_0493_ ), .B2(\LSU/_0476_ ), .ZN(\LSU/_0394_ ) );
OAI21_X1 \LSU/_1051_ ( .A(\LSU/_0471_ ), .B1(\LSU/_0469_ ), .B2(\LSU/_0146_ ), .ZN(\LSU/_0496_ ) );
NOR2_X1 \LSU/_1052_ ( .A1(fanout_net_19 ), .A2(\LSU/_0154_ ), .ZN(\LSU/_0497_ ) );
OAI22_X1 \LSU/_1053_ ( .A1(\LSU/_0496_ ), .A2(\LSU/_0497_ ), .B1(\LSU/_0493_ ), .B2(\LSU/_0477_ ), .ZN(\LSU/_0395_ ) );
OAI21_X1 \LSU/_1054_ ( .A(\LSU/_0471_ ), .B1(\LSU/_0469_ ), .B2(\LSU/_0147_ ), .ZN(\LSU/_0498_ ) );
NOR2_X1 \LSU/_1055_ ( .A1(fanout_net_19 ), .A2(\LSU/_0155_ ), .ZN(\LSU/_0499_ ) );
OAI22_X1 \LSU/_1056_ ( .A1(\LSU/_0498_ ), .A2(\LSU/_0499_ ), .B1(\LSU/_0493_ ), .B2(\LSU/_0478_ ), .ZN(\LSU/_0396_ ) );
OAI21_X1 \LSU/_1057_ ( .A(\LSU/_0471_ ), .B1(\LSU/_0469_ ), .B2(\LSU/_0148_ ), .ZN(\LSU/_0500_ ) );
NOR2_X1 \LSU/_1058_ ( .A1(fanout_net_19 ), .A2(\LSU/_0157_ ), .ZN(\LSU/_0501_ ) );
OAI22_X1 \LSU/_1059_ ( .A1(\LSU/_0500_ ), .A2(\LSU/_0501_ ), .B1(\LSU/_0493_ ), .B2(\LSU/_0479_ ), .ZN(\LSU/_0398_ ) );
OAI21_X1 \LSU/_1060_ ( .A(\LSU/_0471_ ), .B1(\LSU/_0469_ ), .B2(\LSU/_0149_ ), .ZN(\LSU/_0502_ ) );
NOR2_X1 \LSU/_1061_ ( .A1(fanout_net_19 ), .A2(\LSU/_0158_ ), .ZN(\LSU/_0503_ ) );
OAI22_X1 \LSU/_1062_ ( .A1(\LSU/_0502_ ), .A2(\LSU/_0503_ ), .B1(\LSU/_0493_ ), .B2(\LSU/_0480_ ), .ZN(\LSU/_0399_ ) );
OAI21_X1 \LSU/_1063_ ( .A(\LSU/_0471_ ), .B1(\LSU/_0469_ ), .B2(\LSU/_0150_ ), .ZN(\LSU/_0504_ ) );
NOR2_X1 \LSU/_1064_ ( .A1(fanout_net_19 ), .A2(\LSU/_0159_ ), .ZN(\LSU/_0505_ ) );
OAI22_X1 \LSU/_1065_ ( .A1(\LSU/_0504_ ), .A2(\LSU/_0505_ ), .B1(\LSU/_0493_ ), .B2(\LSU/_0481_ ), .ZN(\LSU/_0400_ ) );
OAI21_X1 \LSU/_1066_ ( .A(\LSU/_0471_ ), .B1(\LSU/_0469_ ), .B2(\LSU/_0151_ ), .ZN(\LSU/_0506_ ) );
NOR2_X1 \LSU/_1067_ ( .A1(fanout_net_19 ), .A2(\LSU/_0160_ ), .ZN(\LSU/_0507_ ) );
OAI22_X1 \LSU/_1068_ ( .A1(\LSU/_0506_ ), .A2(\LSU/_0507_ ), .B1(\LSU/_0493_ ), .B2(\LSU/_0482_ ), .ZN(\LSU/_0401_ ) );
MUX2_X1 \LSU/_1069_ ( .A(\LSU/_0161_ ), .B(\LSU/_0152_ ), .S(fanout_net_19 ), .Z(\LSU/_0508_ ) );
MUX2_X1 \LSU/_1070_ ( .A(\LSU/_0508_ ), .B(\LSU/_0483_ ), .S(\LSU/_0327_ ), .Z(\LSU/_0402_ ) );
MUX2_X1 \LSU/_1071_ ( .A(\LSU/_0162_ ), .B(\LSU/_0153_ ), .S(fanout_net_19 ), .Z(\LSU/_0509_ ) );
MUX2_X1 \LSU/_1072_ ( .A(\LSU/_0509_ ), .B(\LSU/_0484_ ), .S(\LSU/_0327_ ), .Z(\LSU/_0403_ ) );
MUX2_X1 \LSU/_1073_ ( .A(\LSU/_0163_ ), .B(\LSU/_0154_ ), .S(fanout_net_19 ), .Z(\LSU/_0510_ ) );
MUX2_X1 \LSU/_1074_ ( .A(\LSU/_0510_ ), .B(\LSU/_0485_ ), .S(\LSU/_0327_ ), .Z(\LSU/_0404_ ) );
MUX2_X1 \LSU/_1075_ ( .A(\LSU/_0164_ ), .B(\LSU/_0155_ ), .S(fanout_net_19 ), .Z(\LSU/_0511_ ) );
MUX2_X1 \LSU/_1076_ ( .A(\LSU/_0511_ ), .B(\LSU/_0486_ ), .S(\LSU/_0327_ ), .Z(\LSU/_0405_ ) );
MUX2_X1 \LSU/_1077_ ( .A(\LSU/_0165_ ), .B(\LSU/_0157_ ), .S(\LSU/_0316_ ), .Z(\LSU/_0512_ ) );
MUX2_X1 \LSU/_1078_ ( .A(\LSU/_0512_ ), .B(\LSU/_0487_ ), .S(\LSU/_0327_ ), .Z(\LSU/_0406_ ) );
MUX2_X1 \LSU/_1079_ ( .A(\LSU/_0166_ ), .B(\LSU/_0158_ ), .S(\LSU/_0316_ ), .Z(\LSU/_0513_ ) );
MUX2_X1 \LSU/_1080_ ( .A(\LSU/_0513_ ), .B(\LSU/_0488_ ), .S(\LSU/_0327_ ), .Z(\LSU/_0407_ ) );
MUX2_X1 \LSU/_1081_ ( .A(\LSU/_0168_ ), .B(\LSU/_0159_ ), .S(\LSU/_0316_ ), .Z(\LSU/_0514_ ) );
MUX2_X1 \LSU/_1082_ ( .A(\LSU/_0514_ ), .B(\LSU/_0489_ ), .S(\LSU/_0327_ ), .Z(\LSU/_0409_ ) );
MUX2_X1 \LSU/_1083_ ( .A(\LSU/_0169_ ), .B(\LSU/_0160_ ), .S(\LSU/_0316_ ), .Z(\LSU/_0515_ ) );
MUX2_X1 \LSU/_1084_ ( .A(\LSU/_0515_ ), .B(\LSU/_0490_ ), .S(\LSU/_0327_ ), .Z(\LSU/_0410_ ) );
INV_X32 \LSU/_1085_ ( .A(\LSU/_0280_ ), .ZN(\LSU/_0516_ ) );
BUF_X32 \LSU/_1086_ ( .A(\LSU/_0516_ ), .Z(\LSU/_0517_ ) );
NAND2_X1 \LSU/_1087_ ( .A1(\LSU/_0517_ ), .A2(\LSU/_0359_ ), .ZN(\LSU/_0518_ ) );
NAND2_X1 \LSU/_1088_ ( .A1(\LSU/_0280_ ), .A2(\LSU/_0368_ ), .ZN(\LSU/_0519_ ) );
NAND2_X1 \LSU/_1089_ ( .A1(\LSU/_0518_ ), .A2(\LSU/_0519_ ), .ZN(\LSU/_0520_ ) );
MUX2_X1 \LSU/_1090_ ( .A(\LSU/_0352_ ), .B(\LSU/_0382_ ), .S(\LSU/_0280_ ), .Z(\LSU/_0521_ ) );
INV_X8 \LSU/_1091_ ( .A(\LSU/_0291_ ), .ZN(\LSU/_0522_ ) );
MUX2_X1 \LSU/_1092_ ( .A(\LSU/_0520_ ), .B(\LSU/_0521_ ), .S(\LSU/_0522_ ), .Z(\LSU/_0523_ ) );
AND2_X4 \LSU/_1093_ ( .A1(\LSU/_0384_ ), .A2(\LSU/_0385_ ), .ZN(\LSU/_0524_ ) );
BUF_X4 \LSU/_1094_ ( .A(\LSU/_0524_ ), .Z(\LSU/_0525_ ) );
BUF_X4 \LSU/_1095_ ( .A(\LSU/_0525_ ), .Z(\LSU/_0526_ ) );
MUX2_X1 \LSU/_1096_ ( .A(\LSU/_0424_ ), .B(\LSU/_0523_ ), .S(\LSU/_0526_ ), .Z(\LSU/_0112_ ) );
NAND2_X1 \LSU/_1097_ ( .A1(\LSU/_0517_ ), .A2(\LSU/_0360_ ), .ZN(\LSU/_0527_ ) );
NAND2_X1 \LSU/_1098_ ( .A1(\LSU/_0280_ ), .A2(\LSU/_0369_ ), .ZN(\LSU/_0528_ ) );
NAND2_X1 \LSU/_1099_ ( .A1(\LSU/_0527_ ), .A2(\LSU/_0528_ ), .ZN(\LSU/_0529_ ) );
MUX2_X1 \LSU/_1100_ ( .A(\LSU/_0363_ ), .B(\LSU/_0383_ ), .S(\LSU/_0280_ ), .Z(\LSU/_0530_ ) );
MUX2_X1 \LSU/_1101_ ( .A(\LSU/_0529_ ), .B(\LSU/_0530_ ), .S(\LSU/_0522_ ), .Z(\LSU/_0531_ ) );
MUX2_X1 \LSU/_1102_ ( .A(\LSU/_0435_ ), .B(\LSU/_0531_ ), .S(\LSU/_0526_ ), .Z(\LSU/_0113_ ) );
NAND2_X1 \LSU/_1103_ ( .A1(\LSU/_0517_ ), .A2(\LSU/_0361_ ), .ZN(\LSU/_0532_ ) );
NAND2_X1 \LSU/_1104_ ( .A1(\LSU/_0280_ ), .A2(\LSU/_0370_ ), .ZN(\LSU/_0533_ ) );
NAND2_X1 \LSU/_1105_ ( .A1(\LSU/_0532_ ), .A2(\LSU/_0533_ ), .ZN(\LSU/_0534_ ) );
MUX2_X1 \LSU/_1106_ ( .A(\LSU/_0374_ ), .B(\LSU/_0353_ ), .S(\LSU/_0280_ ), .Z(\LSU/_0535_ ) );
MUX2_X1 \LSU/_1107_ ( .A(\LSU/_0534_ ), .B(\LSU/_0535_ ), .S(\LSU/_0522_ ), .Z(\LSU/_0536_ ) );
MUX2_X1 \LSU/_1108_ ( .A(\LSU/_0446_ ), .B(\LSU/_0536_ ), .S(\LSU/_0526_ ), .Z(\LSU/_0114_ ) );
NOR2_X1 \LSU/_1109_ ( .A1(\LSU/_0517_ ), .A2(\LSU/_0371_ ), .ZN(\LSU/_0537_ ) );
NOR2_X1 \LSU/_1110_ ( .A1(\LSU/_0280_ ), .A2(\LSU/_0362_ ), .ZN(\LSU/_0538_ ) );
NOR2_X1 \LSU/_1111_ ( .A1(\LSU/_0537_ ), .A2(\LSU/_0538_ ), .ZN(\LSU/_0539_ ) );
MUX2_X1 \LSU/_1112_ ( .A(\LSU/_0377_ ), .B(\LSU/_0354_ ), .S(\LSU/_0280_ ), .Z(\LSU/_0540_ ) );
MUX2_X1 \LSU/_1113_ ( .A(\LSU/_0539_ ), .B(\LSU/_0540_ ), .S(\LSU/_0522_ ), .Z(\LSU/_0541_ ) );
MUX2_X1 \LSU/_1114_ ( .A(\LSU/_0449_ ), .B(\LSU/_0541_ ), .S(\LSU/_0526_ ), .Z(\LSU/_0115_ ) );
NOR2_X1 \LSU/_1115_ ( .A1(\LSU/_0517_ ), .A2(\LSU/_0372_ ), .ZN(\LSU/_0542_ ) );
NOR2_X1 \LSU/_1116_ ( .A1(\LSU/_0280_ ), .A2(\LSU/_0364_ ), .ZN(\LSU/_0543_ ) );
NOR2_X1 \LSU/_1117_ ( .A1(\LSU/_0542_ ), .A2(\LSU/_0543_ ), .ZN(\LSU/_0544_ ) );
MUX2_X1 \LSU/_1118_ ( .A(\LSU/_0378_ ), .B(\LSU/_0355_ ), .S(\LSU/_0280_ ), .Z(\LSU/_0545_ ) );
MUX2_X1 \LSU/_1119_ ( .A(\LSU/_0544_ ), .B(\LSU/_0545_ ), .S(\LSU/_0522_ ), .Z(\LSU/_0546_ ) );
MUX2_X1 \LSU/_1120_ ( .A(\LSU/_0450_ ), .B(\LSU/_0546_ ), .S(\LSU/_0526_ ), .Z(\LSU/_0116_ ) );
NAND2_X1 \LSU/_1121_ ( .A1(\LSU/_0517_ ), .A2(\LSU/_0365_ ), .ZN(\LSU/_0547_ ) );
NAND2_X1 \LSU/_1122_ ( .A1(\LSU/_0280_ ), .A2(\LSU/_0373_ ), .ZN(\LSU/_0548_ ) );
NAND2_X1 \LSU/_1123_ ( .A1(\LSU/_0547_ ), .A2(\LSU/_0548_ ), .ZN(\LSU/_0549_ ) );
MUX2_X1 \LSU/_1124_ ( .A(\LSU/_0379_ ), .B(\LSU/_0356_ ), .S(\LSU/_0280_ ), .Z(\LSU/_0550_ ) );
MUX2_X1 \LSU/_1125_ ( .A(\LSU/_0549_ ), .B(\LSU/_0550_ ), .S(\LSU/_0522_ ), .Z(\LSU/_0551_ ) );
MUX2_X1 \LSU/_1126_ ( .A(\LSU/_0451_ ), .B(\LSU/_0551_ ), .S(\LSU/_0526_ ), .Z(\LSU/_0117_ ) );
NAND2_X1 \LSU/_1127_ ( .A1(\LSU/_0517_ ), .A2(\LSU/_0366_ ), .ZN(\LSU/_0552_ ) );
NAND2_X1 \LSU/_1128_ ( .A1(\LSU/_0280_ ), .A2(\LSU/_0375_ ), .ZN(\LSU/_0553_ ) );
NAND2_X1 \LSU/_1129_ ( .A1(\LSU/_0552_ ), .A2(\LSU/_0553_ ), .ZN(\LSU/_0554_ ) );
MUX2_X1 \LSU/_1130_ ( .A(\LSU/_0380_ ), .B(\LSU/_0357_ ), .S(\LSU/_0280_ ), .Z(\LSU/_0555_ ) );
MUX2_X1 \LSU/_1131_ ( .A(\LSU/_0554_ ), .B(\LSU/_0555_ ), .S(\LSU/_0522_ ), .Z(\LSU/_0556_ ) );
MUX2_X1 \LSU/_1132_ ( .A(\LSU/_0452_ ), .B(\LSU/_0556_ ), .S(\LSU/_0526_ ), .Z(\LSU/_0118_ ) );
AOI21_X1 \LSU/_1133_ ( .A(\LSU/_0453_ ), .B1(\LSU/_0384_ ), .B2(\LSU/_0385_ ), .ZN(\LSU/_0557_ ) );
NAND2_X4 \LSU/_1134_ ( .A1(\LSU/_0516_ ), .A2(\LSU/_0381_ ), .ZN(\LSU/_0558_ ) );
INV_X1 \LSU/_1135_ ( .A(\LSU/_0358_ ), .ZN(\LSU/_0559_ ) );
OAI211_X2 \LSU/_1136_ ( .A(\LSU/_0558_ ), .B(\LSU/_0522_ ), .C1(\LSU/_0559_ ), .C2(\LSU/_0516_ ), .ZN(\LSU/_0560_ ) );
NAND2_X2 \LSU/_1137_ ( .A1(\LSU/_0516_ ), .A2(\LSU/_0367_ ), .ZN(\LSU/_0561_ ) );
NAND2_X2 \LSU/_1138_ ( .A1(\LSU/_0280_ ), .A2(\LSU/_0376_ ), .ZN(\LSU/_0562_ ) );
NAND2_X2 \LSU/_1139_ ( .A1(\LSU/_0561_ ), .A2(\LSU/_0562_ ), .ZN(\LSU/_0563_ ) );
OAI21_X2 \LSU/_1140_ ( .A(\LSU/_0560_ ), .B1(\LSU/_0522_ ), .B2(\LSU/_0563_ ), .ZN(\LSU/_0564_ ) );
AOI21_X1 \LSU/_1141_ ( .A(\LSU/_0557_ ), .B1(\LSU/_0526_ ), .B2(\LSU/_0564_ ), .ZN(\LSU/_0119_ ) );
AND2_X4 \LSU/_1142_ ( .A1(\LSU/_0472_ ), .A2(\LSU/_0144_ ), .ZN(\LSU/_0565_ ) );
NAND2_X1 \LSU/_1143_ ( .A1(\LSU/_0517_ ), .A2(\LSU/_0368_ ), .ZN(\LSU/_0566_ ) );
AOI221_X1 \LSU/_1144_ ( .A(\LSU/_0565_ ), .B1(\LSU/_0291_ ), .B2(\LSU/_0566_ ), .C1(\LSU/_0007_ ), .C2(\LSU/_0473_ ), .ZN(\LSU/_0567_ ) );
MUX2_X1 \LSU/_1145_ ( .A(\LSU/_0382_ ), .B(\LSU/_0359_ ), .S(\LSU/_0280_ ), .Z(\LSU/_0568_ ) );
OAI21_X1 \LSU/_1146_ ( .A(\LSU/_0567_ ), .B1(\LSU/_0291_ ), .B2(\LSU/_0568_ ), .ZN(\LSU/_0569_ ) );
AND2_X4 \LSU/_1147_ ( .A1(\LSU/_0472_ ), .A2(\LSU/_0007_ ), .ZN(\LSU/_0570_ ) );
INV_X2 \LSU/_1148_ ( .A(\LSU/_0570_ ), .ZN(\LSU/_0571_ ) );
NOR2_X4 \LSU/_1149_ ( .A1(\LSU/_0564_ ), .A2(\LSU/_0571_ ), .ZN(\LSU/_0572_ ) );
INV_X1 \LSU/_1150_ ( .A(\LSU/_0572_ ), .ZN(\LSU/_0573_ ) );
NAND2_X1 \LSU/_1151_ ( .A1(\LSU/_0569_ ), .A2(\LSU/_0573_ ), .ZN(\LSU/_0574_ ) );
MUX2_X1 \LSU/_1152_ ( .A(\LSU/_0454_ ), .B(\LSU/_0574_ ), .S(\LSU/_0526_ ), .Z(\LSU/_0120_ ) );
NAND2_X1 \LSU/_1153_ ( .A1(\LSU/_0517_ ), .A2(\LSU/_0369_ ), .ZN(\LSU/_0575_ ) );
AOI221_X1 \LSU/_1154_ ( .A(\LSU/_0565_ ), .B1(\LSU/_0291_ ), .B2(\LSU/_0575_ ), .C1(\LSU/_0007_ ), .C2(\LSU/_0473_ ), .ZN(\LSU/_0576_ ) );
MUX2_X1 \LSU/_1155_ ( .A(\LSU/_0383_ ), .B(\LSU/_0360_ ), .S(\LSU/_0280_ ), .Z(\LSU/_0577_ ) );
OAI21_X1 \LSU/_1156_ ( .A(\LSU/_0576_ ), .B1(\LSU/_0291_ ), .B2(\LSU/_0577_ ), .ZN(\LSU/_0578_ ) );
NAND2_X1 \LSU/_1157_ ( .A1(\LSU/_0578_ ), .A2(\LSU/_0573_ ), .ZN(\LSU/_0579_ ) );
MUX2_X1 \LSU/_1158_ ( .A(\LSU/_0455_ ), .B(\LSU/_0579_ ), .S(\LSU/_0526_ ), .Z(\LSU/_0121_ ) );
NAND2_X1 \LSU/_1159_ ( .A1(\LSU/_0516_ ), .A2(\LSU/_0370_ ), .ZN(\LSU/_0580_ ) );
AOI221_X4 \LSU/_1160_ ( .A(\LSU/_0565_ ), .B1(\LSU/_0291_ ), .B2(\LSU/_0580_ ), .C1(\LSU/_0007_ ), .C2(\LSU/_0473_ ), .ZN(\LSU/_0581_ ) );
MUX2_X1 \LSU/_1161_ ( .A(\LSU/_0353_ ), .B(\LSU/_0361_ ), .S(\LSU/_0280_ ), .Z(\LSU/_0582_ ) );
OAI21_X1 \LSU/_1162_ ( .A(\LSU/_0581_ ), .B1(\LSU/_0291_ ), .B2(\LSU/_0582_ ), .ZN(\LSU/_0583_ ) );
NAND2_X1 \LSU/_1163_ ( .A1(\LSU/_0583_ ), .A2(\LSU/_0573_ ), .ZN(\LSU/_0584_ ) );
BUF_X4 \LSU/_1164_ ( .A(\LSU/_0525_ ), .Z(\LSU/_0585_ ) );
MUX2_X1 \LSU/_1165_ ( .A(\LSU/_0425_ ), .B(\LSU/_0584_ ), .S(\LSU/_0585_ ), .Z(\LSU/_0122_ ) );
NAND2_X1 \LSU/_1166_ ( .A1(\LSU/_0516_ ), .A2(\LSU/_0371_ ), .ZN(\LSU/_0586_ ) );
AOI221_X4 \LSU/_1167_ ( .A(\LSU/_0565_ ), .B1(\LSU/_0291_ ), .B2(\LSU/_0586_ ), .C1(\LSU/_0007_ ), .C2(\LSU/_0473_ ), .ZN(\LSU/_0587_ ) );
MUX2_X1 \LSU/_1168_ ( .A(\LSU/_0354_ ), .B(\LSU/_0362_ ), .S(\LSU/_0280_ ), .Z(\LSU/_0588_ ) );
OAI21_X1 \LSU/_1169_ ( .A(\LSU/_0587_ ), .B1(\LSU/_0291_ ), .B2(\LSU/_0588_ ), .ZN(\LSU/_0589_ ) );
NAND2_X1 \LSU/_1170_ ( .A1(\LSU/_0589_ ), .A2(\LSU/_0573_ ), .ZN(\LSU/_0590_ ) );
MUX2_X1 \LSU/_1171_ ( .A(\LSU/_0426_ ), .B(\LSU/_0590_ ), .S(\LSU/_0585_ ), .Z(\LSU/_0123_ ) );
NAND2_X1 \LSU/_1172_ ( .A1(\LSU/_0516_ ), .A2(\LSU/_0372_ ), .ZN(\LSU/_0591_ ) );
AOI221_X4 \LSU/_1173_ ( .A(\LSU/_0565_ ), .B1(\LSU/_0291_ ), .B2(\LSU/_0591_ ), .C1(\LSU/_0007_ ), .C2(\LSU/_0473_ ), .ZN(\LSU/_0592_ ) );
MUX2_X1 \LSU/_1174_ ( .A(\LSU/_0355_ ), .B(\LSU/_0364_ ), .S(\LSU/_0280_ ), .Z(\LSU/_0593_ ) );
OAI21_X1 \LSU/_1175_ ( .A(\LSU/_0592_ ), .B1(\LSU/_0291_ ), .B2(\LSU/_0593_ ), .ZN(\LSU/_0594_ ) );
NAND2_X1 \LSU/_1176_ ( .A1(\LSU/_0594_ ), .A2(\LSU/_0573_ ), .ZN(\LSU/_0595_ ) );
MUX2_X1 \LSU/_1177_ ( .A(\LSU/_0427_ ), .B(\LSU/_0595_ ), .S(\LSU/_0585_ ), .Z(\LSU/_0124_ ) );
NAND2_X1 \LSU/_1178_ ( .A1(\LSU/_0516_ ), .A2(\LSU/_0373_ ), .ZN(\LSU/_0596_ ) );
AOI221_X4 \LSU/_1179_ ( .A(\LSU/_0565_ ), .B1(\LSU/_0291_ ), .B2(\LSU/_0596_ ), .C1(\LSU/_0007_ ), .C2(\LSU/_0473_ ), .ZN(\LSU/_0597_ ) );
MUX2_X1 \LSU/_1180_ ( .A(\LSU/_0356_ ), .B(\LSU/_0365_ ), .S(\LSU/_0280_ ), .Z(\LSU/_0598_ ) );
OAI21_X1 \LSU/_1181_ ( .A(\LSU/_0597_ ), .B1(\LSU/_0291_ ), .B2(\LSU/_0598_ ), .ZN(\LSU/_0599_ ) );
NAND2_X1 \LSU/_1182_ ( .A1(\LSU/_0599_ ), .A2(\LSU/_0573_ ), .ZN(\LSU/_0600_ ) );
MUX2_X1 \LSU/_1183_ ( .A(\LSU/_0428_ ), .B(\LSU/_0600_ ), .S(\LSU/_0585_ ), .Z(\LSU/_0125_ ) );
NAND2_X1 \LSU/_1184_ ( .A1(\LSU/_0516_ ), .A2(\LSU/_0375_ ), .ZN(\LSU/_0601_ ) );
AOI221_X4 \LSU/_1185_ ( .A(\LSU/_0565_ ), .B1(\LSU/_0291_ ), .B2(\LSU/_0601_ ), .C1(\LSU/_0007_ ), .C2(\LSU/_0473_ ), .ZN(\LSU/_0602_ ) );
MUX2_X1 \LSU/_1186_ ( .A(\LSU/_0357_ ), .B(\LSU/_0366_ ), .S(\LSU/_0280_ ), .Z(\LSU/_0603_ ) );
OAI21_X1 \LSU/_1187_ ( .A(\LSU/_0602_ ), .B1(\LSU/_0291_ ), .B2(\LSU/_0603_ ), .ZN(\LSU/_0604_ ) );
NAND2_X1 \LSU/_1188_ ( .A1(\LSU/_0604_ ), .A2(\LSU/_0573_ ), .ZN(\LSU/_0605_ ) );
MUX2_X1 \LSU/_1189_ ( .A(\LSU/_0429_ ), .B(\LSU/_0605_ ), .S(\LSU/_0585_ ), .Z(\LSU/_0126_ ) );
BUF_X4 \LSU/_1190_ ( .A(\LSU/_0570_ ), .Z(\LSU/_0606_ ) );
OR2_X1 \LSU/_1191_ ( .A1(\LSU/_0606_ ), .A2(\LSU/_0565_ ), .ZN(\LSU/_0607_ ) );
AND3_X4 \LSU/_1192_ ( .A1(\LSU/_0517_ ), .A2(\LSU/_0376_ ), .A3(\LSU/_0291_ ), .ZN(\LSU/_0608_ ) );
MUX2_X1 \LSU/_1193_ ( .A(\LSU/_0358_ ), .B(\LSU/_0367_ ), .S(\LSU/_0280_ ), .Z(\LSU/_0609_ ) );
AOI21_X4 \LSU/_1194_ ( .A(\LSU/_0608_ ), .B1(\LSU/_0609_ ), .B2(\LSU/_0522_ ), .ZN(\LSU/_0610_ ) );
OAI21_X1 \LSU/_1195_ ( .A(\LSU/_0573_ ), .B1(\LSU/_0607_ ), .B2(\LSU/_0610_ ), .ZN(\LSU/_0611_ ) );
MUX2_X1 \LSU/_1196_ ( .A(\LSU/_0430_ ), .B(\LSU/_0611_ ), .S(\LSU/_0585_ ), .Z(\LSU/_0127_ ) );
NOR2_X4 \LSU/_1197_ ( .A1(\LSU/_0467_ ), .A2(\LSU/_0314_ ), .ZN(\LSU/_0612_ ) );
NAND2_X1 \LSU/_1198_ ( .A1(\LSU/_0612_ ), .A2(\LSU/_0007_ ), .ZN(\LSU/_0613_ ) );
BUF_X4 \LSU/_1199_ ( .A(\LSU/_0613_ ), .Z(\LSU/_0614_ ) );
BUF_X8 \LSU/_1200_ ( .A(\LSU/_0572_ ), .Z(\LSU/_0615_ ) );
NAND2_X4 \LSU/_1201_ ( .A1(\LSU/_0466_ ), .A2(\LSU/_0144_ ), .ZN(\LSU/_0616_ ) );
NAND2_X4 \LSU/_1202_ ( .A1(\LSU/_0616_ ), .A2(\LSU/_0006_ ), .ZN(\LSU/_0617_ ) );
BUF_X4 \LSU/_1203_ ( .A(\LSU/_0617_ ), .Z(\LSU/_0618_ ) );
AOI221_X2 \LSU/_1204_ ( .A(\LSU/_0618_ ), .B1(\LSU/_0007_ ), .B2(\LSU/_0473_ ), .C1(\LSU/_0518_ ), .C2(\LSU/_0519_ ), .ZN(\LSU/_0619_ ) );
OAI21_X2 \LSU/_1205_ ( .A(\LSU/_0614_ ), .B1(\LSU/_0615_ ), .B2(\LSU/_0619_ ), .ZN(\LSU/_0620_ ) );
BUF_X4 \LSU/_1206_ ( .A(\LSU/_0610_ ), .Z(\LSU/_0621_ ) );
BUF_X4 \LSU/_1207_ ( .A(\LSU/_0613_ ), .Z(\LSU/_0622_ ) );
OAI21_X1 \LSU/_1208_ ( .A(\LSU/_0620_ ), .B1(\LSU/_0621_ ), .B2(\LSU/_0622_ ), .ZN(\LSU/_0623_ ) );
MUX2_X1 \LSU/_1209_ ( .A(\LSU/_0431_ ), .B(\LSU/_0623_ ), .S(\LSU/_0585_ ), .Z(\LSU/_0128_ ) );
AOI221_X2 \LSU/_1210_ ( .A(\LSU/_0617_ ), .B1(\LSU/_0007_ ), .B2(\LSU/_0473_ ), .C1(\LSU/_0527_ ), .C2(\LSU/_0528_ ), .ZN(\LSU/_0624_ ) );
OAI21_X1 \LSU/_1211_ ( .A(\LSU/_0614_ ), .B1(\LSU/_0615_ ), .B2(\LSU/_0624_ ), .ZN(\LSU/_0625_ ) );
OAI21_X1 \LSU/_1212_ ( .A(\LSU/_0625_ ), .B1(\LSU/_0621_ ), .B2(\LSU/_0622_ ), .ZN(\LSU/_0626_ ) );
MUX2_X1 \LSU/_1213_ ( .A(\LSU/_0432_ ), .B(\LSU/_0626_ ), .S(\LSU/_0585_ ), .Z(\LSU/_0129_ ) );
AOI221_X4 \LSU/_1214_ ( .A(\LSU/_0617_ ), .B1(\LSU/_0007_ ), .B2(\LSU/_0472_ ), .C1(\LSU/_0532_ ), .C2(\LSU/_0533_ ), .ZN(\LSU/_0627_ ) );
OAI21_X2 \LSU/_1215_ ( .A(\LSU/_0614_ ), .B1(\LSU/_0615_ ), .B2(\LSU/_0627_ ), .ZN(\LSU/_0628_ ) );
OAI21_X1 \LSU/_1216_ ( .A(\LSU/_0628_ ), .B1(\LSU/_0621_ ), .B2(\LSU/_0622_ ), .ZN(\LSU/_0629_ ) );
MUX2_X1 \LSU/_1217_ ( .A(\LSU/_0433_ ), .B(\LSU/_0629_ ), .S(\LSU/_0585_ ), .Z(\LSU/_0130_ ) );
NOR4_X1 \LSU/_1218_ ( .A1(\LSU/_0606_ ), .A2(\LSU/_0618_ ), .A3(\LSU/_0538_ ), .A4(\LSU/_0537_ ), .ZN(\LSU/_0630_ ) );
OAI21_X1 \LSU/_1219_ ( .A(\LSU/_0614_ ), .B1(\LSU/_0615_ ), .B2(\LSU/_0630_ ), .ZN(\LSU/_0631_ ) );
OAI21_X1 \LSU/_1220_ ( .A(\LSU/_0631_ ), .B1(\LSU/_0621_ ), .B2(\LSU/_0622_ ), .ZN(\LSU/_0632_ ) );
MUX2_X1 \LSU/_1221_ ( .A(\LSU/_0434_ ), .B(\LSU/_0632_ ), .S(\LSU/_0585_ ), .Z(\LSU/_0131_ ) );
BUF_X4 \LSU/_1222_ ( .A(\LSU/_0613_ ), .Z(\LSU/_0633_ ) );
NOR4_X1 \LSU/_1223_ ( .A1(\LSU/_0606_ ), .A2(\LSU/_0618_ ), .A3(\LSU/_0543_ ), .A4(\LSU/_0542_ ), .ZN(\LSU/_0634_ ) );
OAI21_X1 \LSU/_1224_ ( .A(\LSU/_0633_ ), .B1(\LSU/_0615_ ), .B2(\LSU/_0634_ ), .ZN(\LSU/_0635_ ) );
OAI21_X1 \LSU/_1225_ ( .A(\LSU/_0635_ ), .B1(\LSU/_0621_ ), .B2(\LSU/_0622_ ), .ZN(\LSU/_0636_ ) );
BUF_X4 \LSU/_1226_ ( .A(\LSU/_0525_ ), .Z(\LSU/_0637_ ) );
MUX2_X1 \LSU/_1227_ ( .A(\LSU/_0436_ ), .B(\LSU/_0636_ ), .S(\LSU/_0637_ ), .Z(\LSU/_0132_ ) );
AOI221_X4 \LSU/_1228_ ( .A(\LSU/_0617_ ), .B1(\LSU/_0007_ ), .B2(\LSU/_0472_ ), .C1(\LSU/_0547_ ), .C2(\LSU/_0548_ ), .ZN(\LSU/_0638_ ) );
OAI21_X1 \LSU/_1229_ ( .A(\LSU/_0633_ ), .B1(\LSU/_0615_ ), .B2(\LSU/_0638_ ), .ZN(\LSU/_0639_ ) );
OAI21_X1 \LSU/_1230_ ( .A(\LSU/_0639_ ), .B1(\LSU/_0621_ ), .B2(\LSU/_0622_ ), .ZN(\LSU/_0640_ ) );
MUX2_X1 \LSU/_1231_ ( .A(\LSU/_0437_ ), .B(\LSU/_0640_ ), .S(\LSU/_0637_ ), .Z(\LSU/_0133_ ) );
AOI221_X4 \LSU/_1232_ ( .A(\LSU/_0617_ ), .B1(\LSU/_0007_ ), .B2(\LSU/_0472_ ), .C1(\LSU/_0552_ ), .C2(\LSU/_0553_ ), .ZN(\LSU/_0641_ ) );
OAI21_X2 \LSU/_1233_ ( .A(\LSU/_0633_ ), .B1(\LSU/_0615_ ), .B2(\LSU/_0641_ ), .ZN(\LSU/_0642_ ) );
OAI21_X1 \LSU/_1234_ ( .A(\LSU/_0642_ ), .B1(\LSU/_0621_ ), .B2(\LSU/_0622_ ), .ZN(\LSU/_0643_ ) );
MUX2_X1 \LSU/_1235_ ( .A(\LSU/_0438_ ), .B(\LSU/_0643_ ), .S(\LSU/_0637_ ), .Z(\LSU/_0134_ ) );
AOI221_X4 \LSU/_1236_ ( .A(\LSU/_0617_ ), .B1(\LSU/_0007_ ), .B2(\LSU/_0472_ ), .C1(\LSU/_0561_ ), .C2(\LSU/_0562_ ), .ZN(\LSU/_0644_ ) );
OAI21_X1 \LSU/_1237_ ( .A(\LSU/_0633_ ), .B1(\LSU/_0615_ ), .B2(\LSU/_0644_ ), .ZN(\LSU/_0645_ ) );
OAI21_X1 \LSU/_1238_ ( .A(\LSU/_0645_ ), .B1(\LSU/_0621_ ), .B2(\LSU/_0622_ ), .ZN(\LSU/_0646_ ) );
MUX2_X1 \LSU/_1239_ ( .A(\LSU/_0439_ ), .B(\LSU/_0646_ ), .S(\LSU/_0637_ ), .Z(\LSU/_0135_ ) );
NOR3_X1 \LSU/_1240_ ( .A1(\LSU/_0606_ ), .A2(\LSU/_0618_ ), .A3(\LSU/_0566_ ), .ZN(\LSU/_0647_ ) );
OAI21_X1 \LSU/_1241_ ( .A(\LSU/_0633_ ), .B1(\LSU/_0615_ ), .B2(\LSU/_0647_ ), .ZN(\LSU/_0648_ ) );
OAI21_X1 \LSU/_1242_ ( .A(\LSU/_0648_ ), .B1(\LSU/_0621_ ), .B2(\LSU/_0622_ ), .ZN(\LSU/_0649_ ) );
MUX2_X1 \LSU/_1243_ ( .A(\LSU/_0440_ ), .B(\LSU/_0649_ ), .S(\LSU/_0637_ ), .Z(\LSU/_0136_ ) );
NOR3_X1 \LSU/_1244_ ( .A1(\LSU/_0606_ ), .A2(\LSU/_0618_ ), .A3(\LSU/_0575_ ), .ZN(\LSU/_0650_ ) );
OAI21_X2 \LSU/_1245_ ( .A(\LSU/_0633_ ), .B1(\LSU/_0615_ ), .B2(\LSU/_0650_ ), .ZN(\LSU/_0651_ ) );
OAI21_X1 \LSU/_1246_ ( .A(\LSU/_0651_ ), .B1(\LSU/_0621_ ), .B2(\LSU/_0622_ ), .ZN(\LSU/_0652_ ) );
MUX2_X1 \LSU/_1247_ ( .A(\LSU/_0441_ ), .B(\LSU/_0652_ ), .S(\LSU/_0637_ ), .Z(\LSU/_0137_ ) );
NOR3_X1 \LSU/_1248_ ( .A1(\LSU/_0606_ ), .A2(\LSU/_0618_ ), .A3(\LSU/_0580_ ), .ZN(\LSU/_0653_ ) );
OAI21_X1 \LSU/_1249_ ( .A(\LSU/_0633_ ), .B1(\LSU/_0572_ ), .B2(\LSU/_0653_ ), .ZN(\LSU/_0654_ ) );
OAI21_X1 \LSU/_1250_ ( .A(\LSU/_0654_ ), .B1(\LSU/_0610_ ), .B2(\LSU/_0614_ ), .ZN(\LSU/_0655_ ) );
MUX2_X1 \LSU/_1251_ ( .A(\LSU/_0442_ ), .B(\LSU/_0655_ ), .S(\LSU/_0637_ ), .Z(\LSU/_0138_ ) );
NOR3_X1 \LSU/_1252_ ( .A1(\LSU/_0606_ ), .A2(\LSU/_0618_ ), .A3(\LSU/_0586_ ), .ZN(\LSU/_0656_ ) );
OAI21_X1 \LSU/_1253_ ( .A(\LSU/_0633_ ), .B1(\LSU/_0572_ ), .B2(\LSU/_0656_ ), .ZN(\LSU/_0657_ ) );
OAI21_X1 \LSU/_1254_ ( .A(\LSU/_0657_ ), .B1(\LSU/_0610_ ), .B2(\LSU/_0614_ ), .ZN(\LSU/_0658_ ) );
MUX2_X1 \LSU/_1255_ ( .A(\LSU/_0443_ ), .B(\LSU/_0658_ ), .S(\LSU/_0637_ ), .Z(\LSU/_0139_ ) );
NOR3_X1 \LSU/_1256_ ( .A1(\LSU/_0606_ ), .A2(\LSU/_0618_ ), .A3(\LSU/_0591_ ), .ZN(\LSU/_0659_ ) );
OAI21_X1 \LSU/_1257_ ( .A(\LSU/_0633_ ), .B1(\LSU/_0572_ ), .B2(\LSU/_0659_ ), .ZN(\LSU/_0660_ ) );
OAI21_X1 \LSU/_1258_ ( .A(\LSU/_0660_ ), .B1(\LSU/_0610_ ), .B2(\LSU/_0614_ ), .ZN(\LSU/_0661_ ) );
MUX2_X1 \LSU/_1259_ ( .A(\LSU/_0444_ ), .B(\LSU/_0661_ ), .S(\LSU/_0637_ ), .Z(\LSU/_0140_ ) );
NOR3_X1 \LSU/_1260_ ( .A1(\LSU/_0606_ ), .A2(\LSU/_0618_ ), .A3(\LSU/_0596_ ), .ZN(\LSU/_0662_ ) );
OAI21_X1 \LSU/_1261_ ( .A(\LSU/_0633_ ), .B1(\LSU/_0572_ ), .B2(\LSU/_0662_ ), .ZN(\LSU/_0663_ ) );
OAI21_X1 \LSU/_1262_ ( .A(\LSU/_0663_ ), .B1(\LSU/_0610_ ), .B2(\LSU/_0614_ ), .ZN(\LSU/_0664_ ) );
MUX2_X1 \LSU/_1263_ ( .A(\LSU/_0445_ ), .B(\LSU/_0664_ ), .S(\LSU/_0637_ ), .Z(\LSU/_0141_ ) );
NOR3_X1 \LSU/_1264_ ( .A1(\LSU/_0606_ ), .A2(\LSU/_0618_ ), .A3(\LSU/_0601_ ), .ZN(\LSU/_0665_ ) );
OAI21_X1 \LSU/_1265_ ( .A(\LSU/_0613_ ), .B1(\LSU/_0572_ ), .B2(\LSU/_0665_ ), .ZN(\LSU/_0666_ ) );
OAI21_X1 \LSU/_1266_ ( .A(\LSU/_0666_ ), .B1(\LSU/_0610_ ), .B2(\LSU/_0614_ ), .ZN(\LSU/_0667_ ) );
MUX2_X2 \LSU/_1267_ ( .A(\LSU/_0447_ ), .B(\LSU/_0667_ ), .S(\LSU/_0525_ ), .Z(\LSU/_0142_ ) );
NAND3_X1 \LSU/_1268_ ( .A1(\LSU/_0516_ ), .A2(\LSU/_0376_ ), .A3(\LSU/_0006_ ), .ZN(\LSU/_0668_ ) );
AOI211_X2 \LSU/_1269_ ( .A(\LSU/_0668_ ), .B(\LSU/_0565_ ), .C1(\LSU/_0144_ ), .C2(\LSU/_0612_ ), .ZN(\LSU/_0669_ ) );
AND2_X1 \LSU/_1270_ ( .A1(\LSU/_0669_ ), .A2(\LSU/_0571_ ), .ZN(\LSU/_0670_ ) );
OAI21_X1 \LSU/_1271_ ( .A(\LSU/_0613_ ), .B1(\LSU/_0670_ ), .B2(\LSU/_0572_ ), .ZN(\LSU/_0671_ ) );
OAI21_X1 \LSU/_1272_ ( .A(\LSU/_0671_ ), .B1(\LSU/_0610_ ), .B2(\LSU/_0614_ ), .ZN(\LSU/_0672_ ) );
MUX2_X1 \LSU/_1273_ ( .A(\LSU/_0448_ ), .B(\LSU/_0672_ ), .S(\LSU/_0525_ ), .Z(\LSU/_0143_ ) );
AND2_X2 \LSU/_1274_ ( .A1(\LSU/_0278_ ), .A2(\LSU/_0279_ ), .ZN(\LSU/_0673_ ) );
BUF_X8 \LSU/_1275_ ( .A(\LSU/_0673_ ), .Z(\LSU/_0674_ ) );
BUF_X16 \LSU/_1276_ ( .A(\LSU/_0674_ ), .Z(\LSU/_0675_ ) );
BUF_X16 \LSU/_1277_ ( .A(\LSU/_0675_ ), .Z(\LSU/_0676_ ) );
MUX2_X1 \LSU/_1278_ ( .A(\LSU/_0313_ ), .B(\LSU/_0177_ ), .S(\LSU/_0676_ ), .Z(\LSU/_0013_ ) );
MUX2_X1 \LSU/_1279_ ( .A(\LSU/_0314_ ), .B(\LSU/_0178_ ), .S(\LSU/_0676_ ), .Z(\LSU/_0014_ ) );
MUX2_X1 \LSU/_1280_ ( .A(\LSU/_0144_ ), .B(\LSU/_0179_ ), .S(\LSU/_0676_ ), .Z(\LSU/_0015_ ) );
MUX2_X1 \LSU/_1281_ ( .A(\LSU/_0280_ ), .B(\LSU/_0180_ ), .S(\LSU/_0676_ ), .Z(\LSU/_0016_ ) );
MUX2_X1 \LSU/_1282_ ( .A(\LSU/_0291_ ), .B(\LSU/_0191_ ), .S(\LSU/_0676_ ), .Z(\LSU/_0017_ ) );
MUX2_X1 \LSU/_1283_ ( .A(\LSU/_0302_ ), .B(\LSU/_0202_ ), .S(\LSU/_0676_ ), .Z(\LSU/_0018_ ) );
MUX2_X1 \LSU/_1284_ ( .A(\LSU/_0305_ ), .B(\LSU/_0205_ ), .S(\LSU/_0676_ ), .Z(\LSU/_0019_ ) );
MUX2_X1 \LSU/_1285_ ( .A(\LSU/_0306_ ), .B(\LSU/_0206_ ), .S(\LSU/_0676_ ), .Z(\LSU/_0020_ ) );
MUX2_X1 \LSU/_1286_ ( .A(\LSU/_0307_ ), .B(\LSU/_0207_ ), .S(\LSU/_0676_ ), .Z(\LSU/_0021_ ) );
MUX2_X1 \LSU/_1287_ ( .A(\LSU/_0308_ ), .B(\LSU/_0208_ ), .S(\LSU/_0676_ ), .Z(\LSU/_0022_ ) );
BUF_X4 \LSU/_1288_ ( .A(\LSU/_0674_ ), .Z(\LSU/_0677_ ) );
MUX2_X1 \LSU/_1289_ ( .A(\LSU/_0309_ ), .B(\LSU/_0209_ ), .S(\LSU/_0677_ ), .Z(\LSU/_0023_ ) );
MUX2_X1 \LSU/_1290_ ( .A(\LSU/_0310_ ), .B(\LSU/_0210_ ), .S(\LSU/_0677_ ), .Z(\LSU/_0024_ ) );
MUX2_X1 \LSU/_1291_ ( .A(\LSU/_0311_ ), .B(\LSU/_0211_ ), .S(\LSU/_0677_ ), .Z(\LSU/_0025_ ) );
MUX2_X1 \LSU/_1292_ ( .A(\LSU/_0281_ ), .B(\LSU/_0181_ ), .S(\LSU/_0677_ ), .Z(\LSU/_0026_ ) );
MUX2_X1 \LSU/_1293_ ( .A(\LSU/_0282_ ), .B(\LSU/_0182_ ), .S(\LSU/_0677_ ), .Z(\LSU/_0027_ ) );
MUX2_X1 \LSU/_1294_ ( .A(\LSU/_0283_ ), .B(\LSU/_0183_ ), .S(\LSU/_0677_ ), .Z(\LSU/_0028_ ) );
MUX2_X1 \LSU/_1295_ ( .A(\LSU/_0284_ ), .B(\LSU/_0184_ ), .S(\LSU/_0677_ ), .Z(\LSU/_0029_ ) );
MUX2_X1 \LSU/_1296_ ( .A(\LSU/_0285_ ), .B(\LSU/_0185_ ), .S(\LSU/_0677_ ), .Z(\LSU/_0030_ ) );
MUX2_X1 \LSU/_1297_ ( .A(\LSU/_0286_ ), .B(\LSU/_0186_ ), .S(\LSU/_0677_ ), .Z(\LSU/_0031_ ) );
MUX2_X1 \LSU/_1298_ ( .A(\LSU/_0287_ ), .B(\LSU/_0187_ ), .S(\LSU/_0677_ ), .Z(\LSU/_0032_ ) );
BUF_X4 \LSU/_1299_ ( .A(\LSU/_0674_ ), .Z(\LSU/_0678_ ) );
MUX2_X1 \LSU/_1300_ ( .A(\LSU/_0288_ ), .B(\LSU/_0188_ ), .S(\LSU/_0678_ ), .Z(\LSU/_0033_ ) );
MUX2_X1 \LSU/_1301_ ( .A(\LSU/_0289_ ), .B(\LSU/_0189_ ), .S(\LSU/_0678_ ), .Z(\LSU/_0034_ ) );
MUX2_X1 \LSU/_1302_ ( .A(\LSU/_0290_ ), .B(\LSU/_0190_ ), .S(\LSU/_0678_ ), .Z(\LSU/_0035_ ) );
MUX2_X1 \LSU/_1303_ ( .A(\LSU/_0292_ ), .B(\LSU/_0192_ ), .S(\LSU/_0678_ ), .Z(\LSU/_0036_ ) );
MUX2_X1 \LSU/_1304_ ( .A(\LSU/_0293_ ), .B(\LSU/_0193_ ), .S(\LSU/_0678_ ), .Z(\LSU/_0037_ ) );
MUX2_X1 \LSU/_1305_ ( .A(\LSU/_0294_ ), .B(\LSU/_0194_ ), .S(\LSU/_0678_ ), .Z(\LSU/_0038_ ) );
MUX2_X1 \LSU/_1306_ ( .A(\LSU/_0295_ ), .B(\LSU/_0195_ ), .S(\LSU/_0678_ ), .Z(\LSU/_0039_ ) );
MUX2_X1 \LSU/_1307_ ( .A(\LSU/_0296_ ), .B(\LSU/_0196_ ), .S(\LSU/_0678_ ), .Z(\LSU/_0040_ ) );
MUX2_X1 \LSU/_1308_ ( .A(\LSU/_0297_ ), .B(\LSU/_0197_ ), .S(\LSU/_0678_ ), .Z(\LSU/_0041_ ) );
MUX2_X1 \LSU/_1309_ ( .A(\LSU/_0298_ ), .B(\LSU/_0198_ ), .S(\LSU/_0678_ ), .Z(\LSU/_0042_ ) );
BUF_X4 \LSU/_1310_ ( .A(\LSU/_0674_ ), .Z(\LSU/_0679_ ) );
MUX2_X1 \LSU/_1311_ ( .A(\LSU/_0299_ ), .B(\LSU/_0199_ ), .S(\LSU/_0679_ ), .Z(\LSU/_0043_ ) );
MUX2_X1 \LSU/_1312_ ( .A(\LSU/_0300_ ), .B(\LSU/_0200_ ), .S(\LSU/_0679_ ), .Z(\LSU/_0044_ ) );
MUX2_X1 \LSU/_1313_ ( .A(\LSU/_0301_ ), .B(\LSU/_0201_ ), .S(\LSU/_0679_ ), .Z(\LSU/_0045_ ) );
MUX2_X1 \LSU/_1314_ ( .A(\LSU/_0303_ ), .B(\LSU/_0203_ ), .S(\LSU/_0679_ ), .Z(\LSU/_0046_ ) );
MUX2_X1 \LSU/_1315_ ( .A(\LSU/_0304_ ), .B(\LSU/_0204_ ), .S(\LSU/_0679_ ), .Z(\LSU/_0047_ ) );
MUX2_X1 \LSU/_1316_ ( .A(\LSU/_0316_ ), .B(\LSU/_0213_ ), .S(\LSU/_0679_ ), .Z(\LSU/_0048_ ) );
MUX2_X1 \LSU/_1317_ ( .A(\LSU/_0327_ ), .B(\LSU/_0224_ ), .S(\LSU/_0679_ ), .Z(\LSU/_0049_ ) );
MUX2_X1 \LSU/_1318_ ( .A(\LSU/_0338_ ), .B(\LSU/_0235_ ), .S(\LSU/_0679_ ), .Z(\LSU/_0050_ ) );
MUX2_X1 \LSU/_1319_ ( .A(\LSU/_0341_ ), .B(\LSU/_0238_ ), .S(\LSU/_0679_ ), .Z(\LSU/_0051_ ) );
MUX2_X1 \LSU/_1320_ ( .A(\LSU/_0342_ ), .B(\LSU/_0239_ ), .S(\LSU/_0679_ ), .Z(\LSU/_0052_ ) );
BUF_X4 \LSU/_1321_ ( .A(\LSU/_0674_ ), .Z(\LSU/_0680_ ) );
MUX2_X1 \LSU/_1322_ ( .A(\LSU/_0343_ ), .B(\LSU/_0240_ ), .S(\LSU/_0680_ ), .Z(\LSU/_0053_ ) );
MUX2_X1 \LSU/_1323_ ( .A(\LSU/_0344_ ), .B(\LSU/_0241_ ), .S(\LSU/_0680_ ), .Z(\LSU/_0054_ ) );
MUX2_X1 \LSU/_1324_ ( .A(\LSU/_0345_ ), .B(\LSU/_0242_ ), .S(\LSU/_0680_ ), .Z(\LSU/_0055_ ) );
MUX2_X1 \LSU/_1325_ ( .A(\LSU/_0346_ ), .B(\LSU/_0243_ ), .S(\LSU/_0680_ ), .Z(\LSU/_0056_ ) );
MUX2_X1 \LSU/_1326_ ( .A(\LSU/_0347_ ), .B(\LSU/_0244_ ), .S(\LSU/_0680_ ), .Z(\LSU/_0057_ ) );
MUX2_X1 \LSU/_1327_ ( .A(\LSU/_0317_ ), .B(\LSU/_0214_ ), .S(\LSU/_0680_ ), .Z(\LSU/_0058_ ) );
MUX2_X1 \LSU/_1328_ ( .A(\LSU/_0318_ ), .B(\LSU/_0215_ ), .S(\LSU/_0680_ ), .Z(\LSU/_0059_ ) );
MUX2_X1 \LSU/_1329_ ( .A(\LSU/_0319_ ), .B(\LSU/_0216_ ), .S(\LSU/_0680_ ), .Z(\LSU/_0060_ ) );
MUX2_X1 \LSU/_1330_ ( .A(\LSU/_0320_ ), .B(\LSU/_0217_ ), .S(\LSU/_0680_ ), .Z(\LSU/_0061_ ) );
MUX2_X1 \LSU/_1331_ ( .A(\LSU/_0321_ ), .B(\LSU/_0218_ ), .S(\LSU/_0680_ ), .Z(\LSU/_0062_ ) );
BUF_X4 \LSU/_1332_ ( .A(\LSU/_0674_ ), .Z(\LSU/_0681_ ) );
MUX2_X1 \LSU/_1333_ ( .A(\LSU/_0322_ ), .B(\LSU/_0219_ ), .S(\LSU/_0681_ ), .Z(\LSU/_0063_ ) );
MUX2_X1 \LSU/_1334_ ( .A(\LSU/_0323_ ), .B(\LSU/_0220_ ), .S(\LSU/_0681_ ), .Z(\LSU/_0064_ ) );
MUX2_X1 \LSU/_1335_ ( .A(\LSU/_0324_ ), .B(\LSU/_0221_ ), .S(\LSU/_0681_ ), .Z(\LSU/_0065_ ) );
MUX2_X1 \LSU/_1336_ ( .A(\LSU/_0325_ ), .B(\LSU/_0222_ ), .S(\LSU/_0681_ ), .Z(\LSU/_0066_ ) );
MUX2_X1 \LSU/_1337_ ( .A(\LSU/_0326_ ), .B(\LSU/_0223_ ), .S(\LSU/_0681_ ), .Z(\LSU/_0067_ ) );
MUX2_X1 \LSU/_1338_ ( .A(\LSU/_0328_ ), .B(\LSU/_0225_ ), .S(\LSU/_0681_ ), .Z(\LSU/_0068_ ) );
MUX2_X1 \LSU/_1339_ ( .A(\LSU/_0329_ ), .B(\LSU/_0226_ ), .S(\LSU/_0681_ ), .Z(\LSU/_0069_ ) );
MUX2_X1 \LSU/_1340_ ( .A(\LSU/_0330_ ), .B(\LSU/_0227_ ), .S(\LSU/_0681_ ), .Z(\LSU/_0070_ ) );
MUX2_X1 \LSU/_1341_ ( .A(\LSU/_0331_ ), .B(\LSU/_0228_ ), .S(\LSU/_0681_ ), .Z(\LSU/_0071_ ) );
MUX2_X1 \LSU/_1342_ ( .A(\LSU/_0332_ ), .B(\LSU/_0229_ ), .S(\LSU/_0681_ ), .Z(\LSU/_0072_ ) );
BUF_X4 \LSU/_1343_ ( .A(\LSU/_0674_ ), .Z(\LSU/_0682_ ) );
MUX2_X1 \LSU/_1344_ ( .A(\LSU/_0333_ ), .B(\LSU/_0230_ ), .S(\LSU/_0682_ ), .Z(\LSU/_0073_ ) );
MUX2_X1 \LSU/_1345_ ( .A(\LSU/_0334_ ), .B(\LSU/_0231_ ), .S(\LSU/_0682_ ), .Z(\LSU/_0074_ ) );
MUX2_X1 \LSU/_1346_ ( .A(\LSU/_0335_ ), .B(\LSU/_0232_ ), .S(\LSU/_0682_ ), .Z(\LSU/_0075_ ) );
MUX2_X1 \LSU/_1347_ ( .A(\LSU/_0336_ ), .B(\LSU/_0233_ ), .S(\LSU/_0682_ ), .Z(\LSU/_0076_ ) );
MUX2_X1 \LSU/_1348_ ( .A(\LSU/_0337_ ), .B(\LSU/_0234_ ), .S(\LSU/_0682_ ), .Z(\LSU/_0077_ ) );
MUX2_X1 \LSU/_1349_ ( .A(\LSU/_0339_ ), .B(\LSU/_0236_ ), .S(\LSU/_0682_ ), .Z(\LSU/_0078_ ) );
MUX2_X1 \LSU/_1350_ ( .A(\LSU/_0340_ ), .B(\LSU/_0237_ ), .S(\LSU/_0682_ ), .Z(\LSU/_0079_ ) );
MUX2_X1 \LSU/_1351_ ( .A(\LSU/_0145_ ), .B(\LSU/_0245_ ), .S(\LSU/_0682_ ), .Z(\LSU/_0080_ ) );
MUX2_X1 \LSU/_1352_ ( .A(\LSU/_0156_ ), .B(\LSU/_0256_ ), .S(\LSU/_0682_ ), .Z(\LSU/_0081_ ) );
MUX2_X1 \LSU/_1353_ ( .A(\LSU/_0167_ ), .B(\LSU/_0267_ ), .S(\LSU/_0682_ ), .Z(\LSU/_0082_ ) );
BUF_X4 \LSU/_1354_ ( .A(\LSU/_0674_ ), .Z(\LSU/_0683_ ) );
MUX2_X1 \LSU/_1355_ ( .A(\LSU/_0170_ ), .B(\LSU/_0270_ ), .S(\LSU/_0683_ ), .Z(\LSU/_0083_ ) );
MUX2_X1 \LSU/_1356_ ( .A(\LSU/_0171_ ), .B(\LSU/_0271_ ), .S(\LSU/_0683_ ), .Z(\LSU/_0084_ ) );
MUX2_X1 \LSU/_1357_ ( .A(\LSU/_0172_ ), .B(\LSU/_0272_ ), .S(\LSU/_0683_ ), .Z(\LSU/_0085_ ) );
MUX2_X1 \LSU/_1358_ ( .A(\LSU/_0173_ ), .B(\LSU/_0273_ ), .S(\LSU/_0683_ ), .Z(\LSU/_0086_ ) );
MUX2_X1 \LSU/_1359_ ( .A(\LSU/_0174_ ), .B(\LSU/_0274_ ), .S(\LSU/_0683_ ), .Z(\LSU/_0087_ ) );
MUX2_X1 \LSU/_1360_ ( .A(\LSU/_0175_ ), .B(\LSU/_0275_ ), .S(\LSU/_0683_ ), .Z(\LSU/_0088_ ) );
MUX2_X1 \LSU/_1361_ ( .A(\LSU/_0176_ ), .B(\LSU/_0276_ ), .S(\LSU/_0683_ ), .Z(\LSU/_0089_ ) );
MUX2_X1 \LSU/_1362_ ( .A(\LSU/_0146_ ), .B(\LSU/_0246_ ), .S(\LSU/_0683_ ), .Z(\LSU/_0090_ ) );
MUX2_X1 \LSU/_1363_ ( .A(\LSU/_0147_ ), .B(\LSU/_0247_ ), .S(\LSU/_0683_ ), .Z(\LSU/_0091_ ) );
MUX2_X1 \LSU/_1364_ ( .A(\LSU/_0148_ ), .B(\LSU/_0248_ ), .S(\LSU/_0683_ ), .Z(\LSU/_0092_ ) );
BUF_X4 \LSU/_1365_ ( .A(\LSU/_0674_ ), .Z(\LSU/_0684_ ) );
MUX2_X1 \LSU/_1366_ ( .A(\LSU/_0149_ ), .B(\LSU/_0249_ ), .S(\LSU/_0684_ ), .Z(\LSU/_0093_ ) );
MUX2_X1 \LSU/_1367_ ( .A(\LSU/_0150_ ), .B(\LSU/_0250_ ), .S(\LSU/_0684_ ), .Z(\LSU/_0094_ ) );
MUX2_X1 \LSU/_1368_ ( .A(\LSU/_0151_ ), .B(\LSU/_0251_ ), .S(\LSU/_0684_ ), .Z(\LSU/_0095_ ) );
MUX2_X1 \LSU/_1369_ ( .A(\LSU/_0152_ ), .B(\LSU/_0252_ ), .S(\LSU/_0684_ ), .Z(\LSU/_0096_ ) );
MUX2_X1 \LSU/_1370_ ( .A(\LSU/_0153_ ), .B(\LSU/_0253_ ), .S(\LSU/_0684_ ), .Z(\LSU/_0097_ ) );
MUX2_X1 \LSU/_1371_ ( .A(\LSU/_0154_ ), .B(\LSU/_0254_ ), .S(\LSU/_0684_ ), .Z(\LSU/_0098_ ) );
MUX2_X1 \LSU/_1372_ ( .A(\LSU/_0155_ ), .B(\LSU/_0255_ ), .S(\LSU/_0684_ ), .Z(\LSU/_0099_ ) );
MUX2_X1 \LSU/_1373_ ( .A(\LSU/_0157_ ), .B(\LSU/_0257_ ), .S(\LSU/_0684_ ), .Z(\LSU/_0100_ ) );
MUX2_X1 \LSU/_1374_ ( .A(\LSU/_0158_ ), .B(\LSU/_0258_ ), .S(\LSU/_0684_ ), .Z(\LSU/_0101_ ) );
MUX2_X1 \LSU/_1375_ ( .A(\LSU/_0159_ ), .B(\LSU/_0259_ ), .S(\LSU/_0684_ ), .Z(\LSU/_0102_ ) );
MUX2_X1 \LSU/_1376_ ( .A(\LSU/_0160_ ), .B(\LSU/_0260_ ), .S(\LSU/_0675_ ), .Z(\LSU/_0103_ ) );
MUX2_X1 \LSU/_1377_ ( .A(\LSU/_0161_ ), .B(\LSU/_0261_ ), .S(\LSU/_0675_ ), .Z(\LSU/_0104_ ) );
MUX2_X1 \LSU/_1378_ ( .A(\LSU/_0162_ ), .B(\LSU/_0262_ ), .S(\LSU/_0675_ ), .Z(\LSU/_0105_ ) );
MUX2_X1 \LSU/_1379_ ( .A(\LSU/_0163_ ), .B(\LSU/_0263_ ), .S(\LSU/_0675_ ), .Z(\LSU/_0106_ ) );
MUX2_X1 \LSU/_1380_ ( .A(\LSU/_0164_ ), .B(\LSU/_0264_ ), .S(\LSU/_0675_ ), .Z(\LSU/_0107_ ) );
MUX2_X1 \LSU/_1381_ ( .A(\LSU/_0165_ ), .B(\LSU/_0265_ ), .S(\LSU/_0675_ ), .Z(\LSU/_0108_ ) );
MUX2_X1 \LSU/_1382_ ( .A(\LSU/_0166_ ), .B(\LSU/_0266_ ), .S(\LSU/_0675_ ), .Z(\LSU/_0109_ ) );
MUX2_X1 \LSU/_1383_ ( .A(\LSU/_0168_ ), .B(\LSU/_0268_ ), .S(\LSU/_0675_ ), .Z(\LSU/_0110_ ) );
MUX2_X1 \LSU/_1384_ ( .A(\LSU/_0169_ ), .B(\LSU/_0269_ ), .S(\LSU/_0675_ ), .Z(\LSU/_0111_ ) );
NAND2_X1 \LSU/_1385_ ( .A1(\LSU/_0674_ ), .A2(\LSU/_0212_ ), .ZN(\LSU/_0685_ ) );
INV_X1 \LSU/_1386_ ( .A(\LSU/_0312_ ), .ZN(\LSU/_0686_ ) );
AOI21_X1 \LSU/_1387_ ( .A(\LSU/_0525_ ), .B1(\LSU/_0686_ ), .B2(\LSU/_0315_ ), .ZN(\LSU/_0687_ ) );
NAND3_X1 \LSU/_1388_ ( .A1(\LSU/_0278_ ), .A2(\LSU/_0279_ ), .A3(\LSU/_0277_ ), .ZN(\LSU/_0688_ ) );
AND2_X1 \LSU/_1389_ ( .A1(\LSU/_0418_ ), .A2(\LSU/_0419_ ), .ZN(\LSU/_0689_ ) );
INV_X1 \LSU/_1390_ ( .A(\LSU/_0689_ ), .ZN(\LSU/_0690_ ) );
AND2_X1 \LSU/_1391_ ( .A1(\LSU/_0463_ ), .A2(\LSU/_0459_ ), .ZN(\LSU/_0691_ ) );
NAND2_X1 \LSU/_1392_ ( .A1(\LSU/_0690_ ), .A2(\LSU/_0691_ ), .ZN(\LSU/_0692_ ) );
AND4_X2 \LSU/_1393_ ( .A1(\LSU/_0685_ ), .A2(\LSU/_0687_ ), .A3(\LSU/_0688_ ), .A4(\LSU/_0692_ ), .ZN(\LSU/_0693_ ) );
NOR2_X1 \LSU/_1394_ ( .A1(\LSU/_0461_ ), .A2(\LSU/_0718_ ), .ZN(\LSU/_0694_ ) );
NOR3_X1 \LSU/_1395_ ( .A1(\LSU/_0694_ ), .A2(\LSU/_0460_ ), .A3(\LSU/_0005_ ), .ZN(\LSU/_0695_ ) );
NAND4_X1 \LSU/_1396_ ( .A1(\LSU/_0458_ ), .A2(\LSU/_0718_ ), .A3(\LSU/_0717_ ), .A4(\LSU/_0456_ ), .ZN(\LSU/_0696_ ) );
AND2_X1 \LSU/_1397_ ( .A1(\LSU/_0695_ ), .A2(\LSU/_0696_ ), .ZN(\LSU/_0697_ ) );
INV_X1 \LSU/_1398_ ( .A(\LSU/_0697_ ), .ZN(\LSU/_0698_ ) );
AND3_X1 \LSU/_1399_ ( .A1(\LSU/_0694_ ), .A2(\LSU/_0465_ ), .A3(\LSU/_0351_ ), .ZN(\LSU/_0699_ ) );
AND3_X1 \LSU/_1400_ ( .A1(\LSU/_0718_ ), .A2(\LSU/_0717_ ), .A3(\LSU/_0005_ ), .ZN(\LSU/_0700_ ) );
AOI21_X1 \LSU/_1401_ ( .A(\LSU/_0699_ ), .B1(\LSU/_0690_ ), .B2(\LSU/_0700_ ), .ZN(\LSU/_0701_ ) );
AND2_X1 \LSU/_1402_ ( .A1(\LSU/_0698_ ), .A2(\LSU/_0701_ ), .ZN(\LSU/_0702_ ) );
AOI21_X1 \LSU/_1403_ ( .A(\LSU/_0716_ ), .B1(\LSU/_0693_ ), .B2(\LSU/_0702_ ), .ZN(\LSU/_0010_ ) );
INV_X1 \LSU/_1404_ ( .A(\LSU/_0384_ ), .ZN(\LSU/_0703_ ) );
NAND3_X1 \LSU/_1405_ ( .A1(\LSU/_0694_ ), .A2(\LSU/_0717_ ), .A3(\LSU/_0312_ ), .ZN(\LSU/_0704_ ) );
OR3_X1 \LSU/_1406_ ( .A1(\LSU/_0459_ ), .A2(\LSU/_0717_ ), .A3(\LSU/_0348_ ), .ZN(\LSU/_0705_ ) );
AND4_X1 \LSU/_1407_ ( .A1(\LSU/_0703_ ), .A2(\LSU/_0702_ ), .A3(\LSU/_0704_ ), .A4(\LSU/_0705_ ), .ZN(\LSU/_0706_ ) );
NAND4_X1 \LSU/_1408_ ( .A1(\LSU/_0461_ ), .A2(\LSU/_0717_ ), .A3(\LSU/_0419_ ), .A4(\LSU/_0348_ ), .ZN(\LSU/_0707_ ) );
NOR2_X1 \LSU/_1409_ ( .A1(\LSU/_0464_ ), .A2(\LSU/_0707_ ), .ZN(\LSU/_0708_ ) );
OAI21_X1 \LSU/_1410_ ( .A(\LSU/_0691_ ), .B1(\LSU/_0689_ ), .B2(\LSU/_0348_ ), .ZN(\LSU/_0709_ ) );
OR2_X1 \LSU/_1411_ ( .A1(\LSU/_0708_ ), .A2(\LSU/_0709_ ), .ZN(\LSU/_0710_ ) );
AOI21_X1 \LSU/_1412_ ( .A(\LSU/_0716_ ), .B1(\LSU/_0706_ ), .B2(\LSU/_0710_ ), .ZN(\LSU/_0011_ ) );
NAND4_X1 \LSU/_1413_ ( .A1(\LSU/_0465_ ), .A2(\LSU/_0461_ ), .A3(\LSU/_0718_ ), .A4(\LSU/_0348_ ), .ZN(\LSU/_0711_ ) );
OAI221_X1 \LSU/_1414_ ( .A(\LSU/_0711_ ), .B1(\LSU/_0464_ ), .B2(\LSU/_0707_ ), .C1(\LSU/_0685_ ), .C2(\LSU/_0277_ ), .ZN(\LSU/_0712_ ) );
AND3_X1 \LSU/_1415_ ( .A1(\LSU/_0700_ ), .A2(\LSU/_0418_ ), .A3(\LSU/_0419_ ), .ZN(\LSU/_0713_ ) );
OR2_X1 \LSU/_1416_ ( .A1(\LSU/_0713_ ), .A2(\LSU/_0350_ ), .ZN(\LSU/_0714_ ) );
NOR4_X1 \LSU/_1417_ ( .A1(\LSU/_0712_ ), .A2(\LSU/_0315_ ), .A3(\LSU/_0384_ ), .A4(\LSU/_0714_ ), .ZN(\LSU/_0715_ ) );
AOI21_X1 \LSU/_1418_ ( .A(\LSU/_0716_ ), .B1(\LSU/_0715_ ), .B2(\LSU/_0698_ ), .ZN(\LSU/_0012_ ) );
DFF_X1 \LSU/_1419_ ( .D(\LSU/_0850_ ), .CK(clock ), .Q(\LSU/state [0] ), .QN(\LSU/_0848_ ) );
DFF_X1 \LSU/_1420_ ( .D(\LSU/_0851_ ), .CK(clock ), .Q(\LSU/state [1] ), .QN(\LSU/_0847_ ) );
DFF_X1 \LSU/_1421_ ( .D(\LSU/_0852_ ), .CK(clock ), .Q(\LSU/state [2] ), .QN(\LSU/_0000_ ) );
DFF_X1 \LSU/_1422_ ( .D(\LSU/_0853_ ), .CK(clock ), .Q(\_LSU_io_master_arsize [0] ), .QN(\LSU/_0846_ ) );
DFF_X1 \LSU/_1423_ ( .D(\LSU/_0854_ ), .CK(clock ), .Q(\_LSU_io_master_arsize [1] ), .QN(\LSU/_0845_ ) );
DFF_X1 \LSU/_1424_ ( .D(\LSU/_0855_ ), .CK(clock ), .Q(\LSU/in_memOp [2] ), .QN(\LSU/_0002_ ) );
DFF_X1 \LSU/_1425_ ( .D(\LSU/_0856_ ), .CK(clock ), .Q(\_LSU_io_master_araddr [0] ), .QN(\LSU/_0844_ ) );
DFF_X1 \LSU/_1426_ ( .D(\LSU/_0857_ ), .CK(clock ), .Q(\_LSU_io_master_araddr [1] ), .QN(\LSU/_0001_ ) );
DFF_X1 \LSU/_1427_ ( .D(\LSU/_0858_ ), .CK(clock ), .Q(\_LSU_io_master_araddr [2] ), .QN(\LSU/_0843_ ) );
DFF_X1 \LSU/_1428_ ( .D(\LSU/_0859_ ), .CK(clock ), .Q(\_LSU_io_master_araddr [3] ), .QN(\LSU/_0842_ ) );
DFF_X1 \LSU/_1429_ ( .D(\LSU/_0860_ ), .CK(clock ), .Q(\_LSU_io_master_araddr [4] ), .QN(\LSU/_0841_ ) );
DFF_X1 \LSU/_1430_ ( .D(\LSU/_0861_ ), .CK(clock ), .Q(\_LSU_io_master_araddr [5] ), .QN(\LSU/_0840_ ) );
DFF_X1 \LSU/_1431_ ( .D(\LSU/_0862_ ), .CK(clock ), .Q(\_LSU_io_master_araddr [6] ), .QN(\LSU/_0839_ ) );
DFF_X1 \LSU/_1432_ ( .D(\LSU/_0863_ ), .CK(clock ), .Q(\_LSU_io_master_araddr [7] ), .QN(\LSU/_0838_ ) );
DFF_X1 \LSU/_1433_ ( .D(\LSU/_0864_ ), .CK(clock ), .Q(\_LSU_io_master_araddr [8] ), .QN(\LSU/_0837_ ) );
DFF_X1 \LSU/_1434_ ( .D(\LSU/_0865_ ), .CK(clock ), .Q(\_LSU_io_master_araddr [9] ), .QN(\LSU/_0836_ ) );
DFF_X1 \LSU/_1435_ ( .D(\LSU/_0866_ ), .CK(clock ), .Q(\_LSU_io_master_araddr [10] ), .QN(\LSU/_0835_ ) );
DFF_X1 \LSU/_1436_ ( .D(\LSU/_0867_ ), .CK(clock ), .Q(\_LSU_io_master_araddr [11] ), .QN(\LSU/_0834_ ) );
DFF_X1 \LSU/_1437_ ( .D(\LSU/_0868_ ), .CK(clock ), .Q(\_LSU_io_master_araddr [12] ), .QN(\LSU/_0833_ ) );
DFF_X1 \LSU/_1438_ ( .D(\LSU/_0869_ ), .CK(clock ), .Q(\_LSU_io_master_araddr [13] ), .QN(\LSU/_0832_ ) );
DFF_X1 \LSU/_1439_ ( .D(\LSU/_0870_ ), .CK(clock ), .Q(\_LSU_io_master_araddr [14] ), .QN(\LSU/_0831_ ) );
DFF_X1 \LSU/_1440_ ( .D(\LSU/_0871_ ), .CK(clock ), .Q(\_LSU_io_master_araddr [15] ), .QN(\LSU/_0830_ ) );
DFF_X1 \LSU/_1441_ ( .D(\LSU/_0872_ ), .CK(clock ), .Q(\_LSU_io_master_araddr [16] ), .QN(\LSU/_0829_ ) );
DFF_X1 \LSU/_1442_ ( .D(\LSU/_0873_ ), .CK(clock ), .Q(\_LSU_io_master_araddr [17] ), .QN(\LSU/_0828_ ) );
DFF_X1 \LSU/_1443_ ( .D(\LSU/_0874_ ), .CK(clock ), .Q(\_LSU_io_master_araddr [18] ), .QN(\LSU/_0827_ ) );
DFF_X1 \LSU/_1444_ ( .D(\LSU/_0875_ ), .CK(clock ), .Q(\_LSU_io_master_araddr [19] ), .QN(\LSU/_0826_ ) );
DFF_X1 \LSU/_1445_ ( .D(\LSU/_0876_ ), .CK(clock ), .Q(\_LSU_io_master_araddr [20] ), .QN(\LSU/_0825_ ) );
DFF_X1 \LSU/_1446_ ( .D(\LSU/_0877_ ), .CK(clock ), .Q(\_LSU_io_master_araddr [21] ), .QN(\LSU/_0824_ ) );
DFF_X1 \LSU/_1447_ ( .D(\LSU/_0878_ ), .CK(clock ), .Q(\_LSU_io_master_araddr [22] ), .QN(\LSU/_0823_ ) );
DFF_X1 \LSU/_1448_ ( .D(\LSU/_0879_ ), .CK(clock ), .Q(\_LSU_io_master_araddr [23] ), .QN(\LSU/_0822_ ) );
DFF_X1 \LSU/_1449_ ( .D(\LSU/_0880_ ), .CK(clock ), .Q(\_LSU_io_master_araddr [24] ), .QN(\LSU/_0821_ ) );
DFF_X1 \LSU/_1450_ ( .D(\LSU/_0881_ ), .CK(clock ), .Q(\_LSU_io_master_araddr [25] ), .QN(\LSU/_0820_ ) );
DFF_X1 \LSU/_1451_ ( .D(\LSU/_0882_ ), .CK(clock ), .Q(\_LSU_io_master_araddr [26] ), .QN(\LSU/_0819_ ) );
DFF_X1 \LSU/_1452_ ( .D(\LSU/_0883_ ), .CK(clock ), .Q(\_LSU_io_master_araddr [27] ), .QN(\LSU/_0818_ ) );
DFF_X1 \LSU/_1453_ ( .D(\LSU/_0884_ ), .CK(clock ), .Q(\_LSU_io_master_araddr [28] ), .QN(\LSU/_0817_ ) );
DFF_X1 \LSU/_1454_ ( .D(\LSU/_0885_ ), .CK(clock ), .Q(\_LSU_io_master_araddr [29] ), .QN(\LSU/_0816_ ) );
DFF_X1 \LSU/_1455_ ( .D(\LSU/_0886_ ), .CK(clock ), .Q(\_LSU_io_master_araddr [30] ), .QN(\LSU/_0815_ ) );
DFF_X1 \LSU/_1456_ ( .D(\LSU/_0887_ ), .CK(clock ), .Q(\_LSU_io_master_araddr [31] ), .QN(\LSU/_0814_ ) );
DFF_X1 \LSU/_1457_ ( .D(\LSU/_0888_ ), .CK(clock ), .Q(\_LSU_io_master_awaddr [0] ), .QN(\LSU/_0004_ ) );
DFF_X1 \LSU/_1458_ ( .D(\LSU/_0889_ ), .CK(clock ), .Q(\_LSU_io_master_awaddr [1] ), .QN(\LSU/_0003_ ) );
DFF_X1 \LSU/_1459_ ( .D(\LSU/_0890_ ), .CK(clock ), .Q(\_LSU_io_master_awaddr [2] ), .QN(\LSU/_0813_ ) );
DFF_X1 \LSU/_1460_ ( .D(\LSU/_0891_ ), .CK(clock ), .Q(\_LSU_io_master_awaddr [3] ), .QN(\LSU/_0812_ ) );
DFF_X1 \LSU/_1461_ ( .D(\LSU/_0892_ ), .CK(clock ), .Q(\_LSU_io_master_awaddr [4] ), .QN(\LSU/_0811_ ) );
DFF_X1 \LSU/_1462_ ( .D(\LSU/_0893_ ), .CK(clock ), .Q(\_LSU_io_master_awaddr [5] ), .QN(\LSU/_0810_ ) );
DFF_X1 \LSU/_1463_ ( .D(\LSU/_0894_ ), .CK(clock ), .Q(\_LSU_io_master_awaddr [6] ), .QN(\LSU/_0809_ ) );
DFF_X1 \LSU/_1464_ ( .D(\LSU/_0895_ ), .CK(clock ), .Q(\_LSU_io_master_awaddr [7] ), .QN(\LSU/_0808_ ) );
DFF_X1 \LSU/_1465_ ( .D(\LSU/_0896_ ), .CK(clock ), .Q(\_LSU_io_master_awaddr [8] ), .QN(\LSU/_0807_ ) );
DFF_X1 \LSU/_1466_ ( .D(\LSU/_0897_ ), .CK(clock ), .Q(\_LSU_io_master_awaddr [9] ), .QN(\LSU/_0806_ ) );
DFF_X1 \LSU/_1467_ ( .D(\LSU/_0898_ ), .CK(clock ), .Q(\_LSU_io_master_awaddr [10] ), .QN(\LSU/_0805_ ) );
DFF_X1 \LSU/_1468_ ( .D(\LSU/_0899_ ), .CK(clock ), .Q(\_LSU_io_master_awaddr [11] ), .QN(\LSU/_0804_ ) );
DFF_X1 \LSU/_1469_ ( .D(\LSU/_0900_ ), .CK(clock ), .Q(\_LSU_io_master_awaddr [12] ), .QN(\LSU/_0803_ ) );
DFF_X1 \LSU/_1470_ ( .D(\LSU/_0901_ ), .CK(clock ), .Q(\_LSU_io_master_awaddr [13] ), .QN(\LSU/_0802_ ) );
DFF_X1 \LSU/_1471_ ( .D(\LSU/_0902_ ), .CK(clock ), .Q(\_LSU_io_master_awaddr [14] ), .QN(\LSU/_0801_ ) );
DFF_X1 \LSU/_1472_ ( .D(\LSU/_0903_ ), .CK(clock ), .Q(\_LSU_io_master_awaddr [15] ), .QN(\LSU/_0800_ ) );
DFF_X1 \LSU/_1473_ ( .D(\LSU/_0904_ ), .CK(clock ), .Q(\_LSU_io_master_awaddr [16] ), .QN(\LSU/_0799_ ) );
DFF_X1 \LSU/_1474_ ( .D(\LSU/_0905_ ), .CK(clock ), .Q(\_LSU_io_master_awaddr [17] ), .QN(\LSU/_0798_ ) );
DFF_X1 \LSU/_1475_ ( .D(\LSU/_0906_ ), .CK(clock ), .Q(\_LSU_io_master_awaddr [18] ), .QN(\LSU/_0797_ ) );
DFF_X1 \LSU/_1476_ ( .D(\LSU/_0907_ ), .CK(clock ), .Q(\_LSU_io_master_awaddr [19] ), .QN(\LSU/_0796_ ) );
DFF_X1 \LSU/_1477_ ( .D(\LSU/_0908_ ), .CK(clock ), .Q(\_LSU_io_master_awaddr [20] ), .QN(\LSU/_0795_ ) );
DFF_X1 \LSU/_1478_ ( .D(\LSU/_0909_ ), .CK(clock ), .Q(\_LSU_io_master_awaddr [21] ), .QN(\LSU/_0794_ ) );
DFF_X1 \LSU/_1479_ ( .D(\LSU/_0910_ ), .CK(clock ), .Q(\_LSU_io_master_awaddr [22] ), .QN(\LSU/_0793_ ) );
DFF_X1 \LSU/_1480_ ( .D(\LSU/_0911_ ), .CK(clock ), .Q(\_LSU_io_master_awaddr [23] ), .QN(\LSU/_0792_ ) );
DFF_X1 \LSU/_1481_ ( .D(\LSU/_0912_ ), .CK(clock ), .Q(\_LSU_io_master_awaddr [24] ), .QN(\LSU/_0791_ ) );
DFF_X1 \LSU/_1482_ ( .D(\LSU/_0913_ ), .CK(clock ), .Q(\_LSU_io_master_awaddr [25] ), .QN(\LSU/_0790_ ) );
DFF_X1 \LSU/_1483_ ( .D(\LSU/_0914_ ), .CK(clock ), .Q(\_LSU_io_master_awaddr [26] ), .QN(\LSU/_0789_ ) );
DFF_X1 \LSU/_1484_ ( .D(\LSU/_0915_ ), .CK(clock ), .Q(\_LSU_io_master_awaddr [27] ), .QN(\LSU/_0788_ ) );
DFF_X1 \LSU/_1485_ ( .D(\LSU/_0916_ ), .CK(clock ), .Q(\_LSU_io_master_awaddr [28] ), .QN(\LSU/_0787_ ) );
DFF_X1 \LSU/_1486_ ( .D(\LSU/_0917_ ), .CK(clock ), .Q(\_LSU_io_master_awaddr [29] ), .QN(\LSU/_0786_ ) );
DFF_X1 \LSU/_1487_ ( .D(\LSU/_0918_ ), .CK(clock ), .Q(\_LSU_io_master_awaddr [30] ), .QN(\LSU/_0785_ ) );
DFF_X1 \LSU/_1488_ ( .D(\LSU/_0919_ ), .CK(clock ), .Q(\_LSU_io_master_awaddr [31] ), .QN(\LSU/_0784_ ) );
DFF_X1 \LSU/_1489_ ( .D(\LSU/_0920_ ), .CK(clock ), .Q(\LSU/in_wdata [0] ), .QN(\LSU/_0783_ ) );
DFF_X1 \LSU/_1490_ ( .D(\LSU/_0921_ ), .CK(clock ), .Q(\LSU/in_wdata [1] ), .QN(\LSU/_0782_ ) );
DFF_X1 \LSU/_1491_ ( .D(\LSU/_0922_ ), .CK(clock ), .Q(\LSU/in_wdata [2] ), .QN(\LSU/_0781_ ) );
DFF_X1 \LSU/_1492_ ( .D(\LSU/_0923_ ), .CK(clock ), .Q(\LSU/in_wdata [3] ), .QN(\LSU/_0780_ ) );
DFF_X1 \LSU/_1493_ ( .D(\LSU/_0924_ ), .CK(clock ), .Q(\LSU/in_wdata [4] ), .QN(\LSU/_0779_ ) );
DFF_X1 \LSU/_1494_ ( .D(\LSU/_0925_ ), .CK(clock ), .Q(\LSU/in_wdata [5] ), .QN(\LSU/_0778_ ) );
DFF_X1 \LSU/_1495_ ( .D(\LSU/_0926_ ), .CK(clock ), .Q(\LSU/in_wdata [6] ), .QN(\LSU/_0777_ ) );
DFF_X1 \LSU/_1496_ ( .D(\LSU/_0927_ ), .CK(clock ), .Q(\LSU/in_wdata [7] ), .QN(\LSU/_0776_ ) );
DFF_X1 \LSU/_1497_ ( .D(\LSU/_0928_ ), .CK(clock ), .Q(\LSU/in_wdata [8] ), .QN(\LSU/_0775_ ) );
DFF_X1 \LSU/_1498_ ( .D(\LSU/_0929_ ), .CK(clock ), .Q(\LSU/in_wdata [9] ), .QN(\LSU/_0774_ ) );
DFF_X1 \LSU/_1499_ ( .D(\LSU/_0930_ ), .CK(clock ), .Q(\LSU/in_wdata [10] ), .QN(\LSU/_0773_ ) );
DFF_X1 \LSU/_1500_ ( .D(\LSU/_0931_ ), .CK(clock ), .Q(\LSU/in_wdata [11] ), .QN(\LSU/_0772_ ) );
DFF_X1 \LSU/_1501_ ( .D(\LSU/_0932_ ), .CK(clock ), .Q(\LSU/in_wdata [12] ), .QN(\LSU/_0771_ ) );
DFF_X1 \LSU/_1502_ ( .D(\LSU/_0933_ ), .CK(clock ), .Q(\LSU/in_wdata [13] ), .QN(\LSU/_0770_ ) );
DFF_X1 \LSU/_1503_ ( .D(\LSU/_0934_ ), .CK(clock ), .Q(\LSU/in_wdata [14] ), .QN(\LSU/_0769_ ) );
DFF_X1 \LSU/_1504_ ( .D(\LSU/_0935_ ), .CK(clock ), .Q(\LSU/in_wdata [15] ), .QN(\LSU/_0768_ ) );
DFF_X1 \LSU/_1505_ ( .D(\LSU/_0936_ ), .CK(clock ), .Q(\LSU/in_wdata [16] ), .QN(\LSU/_0767_ ) );
DFF_X1 \LSU/_1506_ ( .D(\LSU/_0937_ ), .CK(clock ), .Q(\LSU/in_wdata [17] ), .QN(\LSU/_0766_ ) );
DFF_X1 \LSU/_1507_ ( .D(\LSU/_0938_ ), .CK(clock ), .Q(\LSU/in_wdata [18] ), .QN(\LSU/_0765_ ) );
DFF_X1 \LSU/_1508_ ( .D(\LSU/_0939_ ), .CK(clock ), .Q(\LSU/in_wdata [19] ), .QN(\LSU/_0764_ ) );
DFF_X1 \LSU/_1509_ ( .D(\LSU/_0940_ ), .CK(clock ), .Q(\LSU/in_wdata [20] ), .QN(\LSU/_0763_ ) );
DFF_X1 \LSU/_1510_ ( .D(\LSU/_0941_ ), .CK(clock ), .Q(\LSU/in_wdata [21] ), .QN(\LSU/_0762_ ) );
DFF_X1 \LSU/_1511_ ( .D(\LSU/_0942_ ), .CK(clock ), .Q(\LSU/in_wdata [22] ), .QN(\LSU/_0761_ ) );
DFF_X1 \LSU/_1512_ ( .D(\LSU/_0943_ ), .CK(clock ), .Q(\LSU/in_wdata [23] ), .QN(\LSU/_0760_ ) );
DFF_X1 \LSU/_1513_ ( .D(\LSU/_0944_ ), .CK(clock ), .Q(\LSU/in_wdata [24] ), .QN(\LSU/_0759_ ) );
DFF_X1 \LSU/_1514_ ( .D(\LSU/_0945_ ), .CK(clock ), .Q(\LSU/in_wdata [25] ), .QN(\LSU/_0758_ ) );
DFF_X1 \LSU/_1515_ ( .D(\LSU/_0946_ ), .CK(clock ), .Q(\LSU/in_wdata [26] ), .QN(\LSU/_0757_ ) );
DFF_X1 \LSU/_1516_ ( .D(\LSU/_0947_ ), .CK(clock ), .Q(\LSU/in_wdata [27] ), .QN(\LSU/_0756_ ) );
DFF_X1 \LSU/_1517_ ( .D(\LSU/_0948_ ), .CK(clock ), .Q(\LSU/in_wdata [28] ), .QN(\LSU/_0755_ ) );
DFF_X1 \LSU/_1518_ ( .D(\LSU/_0949_ ), .CK(clock ), .Q(\LSU/in_wdata [29] ), .QN(\LSU/_0754_ ) );
DFF_X1 \LSU/_1519_ ( .D(\LSU/_0950_ ), .CK(clock ), .Q(\LSU/in_wdata [30] ), .QN(\LSU/_0753_ ) );
DFF_X1 \LSU/_1520_ ( .D(\LSU/_0951_ ), .CK(clock ), .Q(\LSU/in_wdata [31] ), .QN(\LSU/_0752_ ) );
DFF_X1 \LSU/_1521_ ( .D(\LSU/_0952_ ), .CK(clock ), .Q(\_LSU_io_out_bits_rdata [0] ), .QN(\LSU/_0751_ ) );
DFF_X1 \LSU/_1522_ ( .D(\LSU/_0953_ ), .CK(clock ), .Q(\_LSU_io_out_bits_rdata [1] ), .QN(\LSU/_0750_ ) );
DFF_X1 \LSU/_1523_ ( .D(\LSU/_0954_ ), .CK(clock ), .Q(\_LSU_io_out_bits_rdata [2] ), .QN(\LSU/_0749_ ) );
DFF_X1 \LSU/_1524_ ( .D(\LSU/_0955_ ), .CK(clock ), .Q(\_LSU_io_out_bits_rdata [3] ), .QN(\LSU/_0748_ ) );
DFF_X1 \LSU/_1525_ ( .D(\LSU/_0956_ ), .CK(clock ), .Q(\_LSU_io_out_bits_rdata [4] ), .QN(\LSU/_0747_ ) );
DFF_X1 \LSU/_1526_ ( .D(\LSU/_0957_ ), .CK(clock ), .Q(\_LSU_io_out_bits_rdata [5] ), .QN(\LSU/_0746_ ) );
DFF_X1 \LSU/_1527_ ( .D(\LSU/_0958_ ), .CK(clock ), .Q(\_LSU_io_out_bits_rdata [6] ), .QN(\LSU/_0745_ ) );
DFF_X1 \LSU/_1528_ ( .D(\LSU/_0959_ ), .CK(clock ), .Q(\_LSU_io_out_bits_rdata [7] ), .QN(\LSU/_0744_ ) );
DFF_X1 \LSU/_1529_ ( .D(\LSU/_0960_ ), .CK(clock ), .Q(\_LSU_io_out_bits_rdata [8] ), .QN(\LSU/_0743_ ) );
DFF_X1 \LSU/_1530_ ( .D(\LSU/_0961_ ), .CK(clock ), .Q(\_LSU_io_out_bits_rdata [9] ), .QN(\LSU/_0742_ ) );
DFF_X1 \LSU/_1531_ ( .D(\LSU/_0962_ ), .CK(clock ), .Q(\_LSU_io_out_bits_rdata [10] ), .QN(\LSU/_0741_ ) );
DFF_X1 \LSU/_1532_ ( .D(\LSU/_0963_ ), .CK(clock ), .Q(\_LSU_io_out_bits_rdata [11] ), .QN(\LSU/_0740_ ) );
DFF_X1 \LSU/_1533_ ( .D(\LSU/_0964_ ), .CK(clock ), .Q(\_LSU_io_out_bits_rdata [12] ), .QN(\LSU/_0739_ ) );
DFF_X1 \LSU/_1534_ ( .D(\LSU/_0965_ ), .CK(clock ), .Q(\_LSU_io_out_bits_rdata [13] ), .QN(\LSU/_0738_ ) );
DFF_X1 \LSU/_1535_ ( .D(\LSU/_0966_ ), .CK(clock ), .Q(\_LSU_io_out_bits_rdata [14] ), .QN(\LSU/_0737_ ) );
DFF_X1 \LSU/_1536_ ( .D(\LSU/_0967_ ), .CK(clock ), .Q(\_LSU_io_out_bits_rdata [15] ), .QN(\LSU/_0736_ ) );
DFF_X1 \LSU/_1537_ ( .D(\LSU/_0968_ ), .CK(clock ), .Q(\_LSU_io_out_bits_rdata [16] ), .QN(\LSU/_0735_ ) );
DFF_X1 \LSU/_1538_ ( .D(\LSU/_0969_ ), .CK(clock ), .Q(\_LSU_io_out_bits_rdata [17] ), .QN(\LSU/_0734_ ) );
DFF_X1 \LSU/_1539_ ( .D(\LSU/_0970_ ), .CK(clock ), .Q(\_LSU_io_out_bits_rdata [18] ), .QN(\LSU/_0733_ ) );
DFF_X1 \LSU/_1540_ ( .D(\LSU/_0971_ ), .CK(clock ), .Q(\_LSU_io_out_bits_rdata [19] ), .QN(\LSU/_0732_ ) );
DFF_X1 \LSU/_1541_ ( .D(\LSU/_0972_ ), .CK(clock ), .Q(\_LSU_io_out_bits_rdata [20] ), .QN(\LSU/_0731_ ) );
DFF_X1 \LSU/_1542_ ( .D(\LSU/_0973_ ), .CK(clock ), .Q(\_LSU_io_out_bits_rdata [21] ), .QN(\LSU/_0730_ ) );
DFF_X1 \LSU/_1543_ ( .D(\LSU/_0974_ ), .CK(clock ), .Q(\_LSU_io_out_bits_rdata [22] ), .QN(\LSU/_0729_ ) );
DFF_X1 \LSU/_1544_ ( .D(\LSU/_0975_ ), .CK(clock ), .Q(\_LSU_io_out_bits_rdata [23] ), .QN(\LSU/_0728_ ) );
DFF_X1 \LSU/_1545_ ( .D(\LSU/_0976_ ), .CK(clock ), .Q(\_LSU_io_out_bits_rdata [24] ), .QN(\LSU/_0727_ ) );
DFF_X1 \LSU/_1546_ ( .D(\LSU/_0977_ ), .CK(clock ), .Q(\_LSU_io_out_bits_rdata [25] ), .QN(\LSU/_0726_ ) );
DFF_X1 \LSU/_1547_ ( .D(\LSU/_0978_ ), .CK(clock ), .Q(\_LSU_io_out_bits_rdata [26] ), .QN(\LSU/_0725_ ) );
DFF_X1 \LSU/_1548_ ( .D(\LSU/_0979_ ), .CK(clock ), .Q(\_LSU_io_out_bits_rdata [27] ), .QN(\LSU/_0724_ ) );
DFF_X1 \LSU/_1549_ ( .D(\LSU/_0980_ ), .CK(clock ), .Q(\_LSU_io_out_bits_rdata [28] ), .QN(\LSU/_0723_ ) );
DFF_X1 \LSU/_1550_ ( .D(\LSU/_0981_ ), .CK(clock ), .Q(\_LSU_io_out_bits_rdata [29] ), .QN(\LSU/_0722_ ) );
DFF_X1 \LSU/_1551_ ( .D(\LSU/_0982_ ), .CK(clock ), .Q(\_LSU_io_out_bits_rdata [30] ), .QN(\LSU/_0721_ ) );
DFF_X1 \LSU/_1552_ ( .D(\LSU/_0983_ ), .CK(clock ), .Q(\_LSU_io_out_bits_rdata [31] ), .QN(\LSU/_0720_ ) );
LOGIC0_X1 \LSU/_1553_ ( .Z(\LSU/_0849_ ) );
BUF_X1 \LSU/_1554_ ( .A(\_LSU_io_master_arsize [0] ), .Z(\LSU/in_memOp [0] ) );
BUF_X1 \LSU/_1555_ ( .A(\_LSU_io_master_arsize [1] ), .Z(\LSU/in_memOp [1] ) );
BUF_X1 \LSU/_1556_ ( .A(\LSU/_0849_ ), .Z(\_LSU_io_master_arsize [2] ) );
BUF_X1 \LSU/_1557_ ( .A(\_LSU_io_master_arsize [0] ), .Z(\_LSU_io_master_awsize [0] ) );
BUF_X1 \LSU/_1558_ ( .A(\_LSU_io_master_arsize [1] ), .Z(\_LSU_io_master_awsize [1] ) );
BUF_X1 \LSU/_1559_ ( .A(\LSU/_0849_ ), .Z(\_LSU_io_master_awsize [2] ) );
BUF_X1 \LSU/_1560_ ( .A(_LSU_io_master_wlast ), .Z(_LSU_io_master_wvalid ) );
BUF_X1 \LSU/_1561_ ( .A(\LSU/state [1] ), .Z(\LSU/_0718_ ) );
BUF_X1 \LSU/_1562_ ( .A(\LSU/state [0] ), .Z(\LSU/_0717_ ) );
BUF_X1 \LSU/_1563_ ( .A(\LSU/_0000_ ), .Z(\LSU/_0005_ ) );
BUF_X1 \LSU/_1564_ ( .A(\LSU/_0457_ ), .Z(_LSU_io_out_valid ) );
BUF_X1 \LSU/_1565_ ( .A(\LSU/state [2] ), .Z(\LSU/_0719_ ) );
BUF_X1 \LSU/_1566_ ( .A(\LSU/_0315_ ), .Z(_LSU_io_master_arvalid ) );
BUF_X1 \LSU/_1567_ ( .A(\LSU/_0384_ ), .Z(_LSU_io_master_rready ) );
BUF_X1 \LSU/_1568_ ( .A(\LSU/_0350_ ), .Z(_LSU_io_master_bready ) );
BUF_X1 \LSU/_1569_ ( .A(\LSU/_0349_ ), .Z(_LSU_io_master_awvalid ) );
BUF_X1 \LSU/_1570_ ( .A(\LSU/_0278_ ), .Z(_LSU_io_in_ready ) );
BUF_X1 \LSU/_1571_ ( .A(_AXI4Interconnect_io_fanIn_1_rvalid ), .Z(\LSU/_0385_ ) );
BUF_X1 \LSU/_1572_ ( .A(\_AXI4Interconnect_io_fanIn_1_rdata [7] ), .Z(\LSU/_0381_ ) );
BUF_X1 \LSU/_1573_ ( .A(\_AXI4Interconnect_io_fanIn_1_rdata [15] ), .Z(\LSU/_0358_ ) );
BUF_X1 \LSU/_1574_ ( .A(\_LSU_io_master_araddr [0] ), .Z(\LSU/_0280_ ) );
BUF_X1 \LSU/_1575_ ( .A(\_AXI4Interconnect_io_fanIn_1_rdata [23] ), .Z(\LSU/_0367_ ) );
BUF_X1 \LSU/_1576_ ( .A(\_AXI4Interconnect_io_fanIn_1_rdata [31] ), .Z(\LSU/_0376_ ) );
BUF_X1 \LSU/_1577_ ( .A(\_LSU_io_master_araddr [1] ), .Z(\LSU/_0291_ ) );
BUF_X1 \LSU/_1578_ ( .A(\_AXI4Interconnect_io_fanIn_1_rdata [8] ), .Z(\LSU/_0382_ ) );
BUF_X1 \LSU/_1579_ ( .A(\_AXI4Interconnect_io_fanIn_1_rdata [16] ), .Z(\LSU/_0359_ ) );
BUF_X1 \LSU/_1580_ ( .A(\_AXI4Interconnect_io_fanIn_1_rdata [24] ), .Z(\LSU/_0368_ ) );
BUF_X1 \LSU/_1581_ ( .A(\_LSU_io_master_arsize [1] ), .Z(\LSU/_0314_ ) );
BUF_X1 \LSU/_1582_ ( .A(\_LSU_io_master_arsize [0] ), .Z(\LSU/_0313_ ) );
BUF_X1 \LSU/_1583_ ( .A(\LSU/_0002_ ), .Z(\LSU/_0007_ ) );
BUF_X1 \LSU/_1584_ ( .A(\LSU/in_memOp [2] ), .Z(\LSU/_0144_ ) );
BUF_X1 \LSU/_1585_ ( .A(\_AXI4Interconnect_io_fanIn_1_rdata [9] ), .Z(\LSU/_0383_ ) );
BUF_X1 \LSU/_1586_ ( .A(\_AXI4Interconnect_io_fanIn_1_rdata [17] ), .Z(\LSU/_0360_ ) );
BUF_X1 \LSU/_1587_ ( .A(\_AXI4Interconnect_io_fanIn_1_rdata [25] ), .Z(\LSU/_0369_ ) );
BUF_X1 \LSU/_1588_ ( .A(\_AXI4Interconnect_io_fanIn_1_rdata [10] ), .Z(\LSU/_0353_ ) );
BUF_X1 \LSU/_1589_ ( .A(\_AXI4Interconnect_io_fanIn_1_rdata [18] ), .Z(\LSU/_0361_ ) );
BUF_X1 \LSU/_1590_ ( .A(\_AXI4Interconnect_io_fanIn_1_rdata [26] ), .Z(\LSU/_0370_ ) );
BUF_X1 \LSU/_1591_ ( .A(\_AXI4Interconnect_io_fanIn_1_rdata [11] ), .Z(\LSU/_0354_ ) );
BUF_X1 \LSU/_1592_ ( .A(\_AXI4Interconnect_io_fanIn_1_rdata [19] ), .Z(\LSU/_0362_ ) );
BUF_X1 \LSU/_1593_ ( .A(\_AXI4Interconnect_io_fanIn_1_rdata [27] ), .Z(\LSU/_0371_ ) );
BUF_X1 \LSU/_1594_ ( .A(\_AXI4Interconnect_io_fanIn_1_rdata [12] ), .Z(\LSU/_0355_ ) );
BUF_X1 \LSU/_1595_ ( .A(\_AXI4Interconnect_io_fanIn_1_rdata [20] ), .Z(\LSU/_0364_ ) );
BUF_X1 \LSU/_1596_ ( .A(\_AXI4Interconnect_io_fanIn_1_rdata [28] ), .Z(\LSU/_0372_ ) );
BUF_X1 \LSU/_1597_ ( .A(\_AXI4Interconnect_io_fanIn_1_rdata [13] ), .Z(\LSU/_0356_ ) );
BUF_X1 \LSU/_1598_ ( .A(\_AXI4Interconnect_io_fanIn_1_rdata [21] ), .Z(\LSU/_0365_ ) );
BUF_X1 \LSU/_1599_ ( .A(\_AXI4Interconnect_io_fanIn_1_rdata [29] ), .Z(\LSU/_0373_ ) );
BUF_X1 \LSU/_1600_ ( .A(\_AXI4Interconnect_io_fanIn_1_rdata [14] ), .Z(\LSU/_0357_ ) );
BUF_X1 \LSU/_1601_ ( .A(\_AXI4Interconnect_io_fanIn_1_rdata [22] ), .Z(\LSU/_0366_ ) );
BUF_X1 \LSU/_1602_ ( .A(\_AXI4Interconnect_io_fanIn_1_rdata [30] ), .Z(\LSU/_0375_ ) );
BUF_X1 \LSU/_1603_ ( .A(\LSU/_0001_ ), .Z(\LSU/_0006_ ) );
BUF_X1 \LSU/_1604_ ( .A(_EXU_io_LSUOut_ready ), .Z(\LSU/_0456_ ) );
BUF_X1 \LSU/_1605_ ( .A(_AXI4Interconnect_io_fanIn_1_arready ), .Z(\LSU/_0312_ ) );
BUF_X1 \LSU/_1606_ ( .A(_AXI4Interconnect_io_fanIn_1_bvalid ), .Z(\LSU/_0351_ ) );
BUF_X1 \LSU/_1607_ ( .A(_AXI4Interconnect_io_fanIn_1_wready ), .Z(\LSU/_0419_ ) );
BUF_X1 \LSU/_1608_ ( .A(_AXI4Interconnect_io_fanIn_1_awready ), .Z(\LSU/_0348_ ) );
BUF_X1 \LSU/_1609_ ( .A(_EXU_io_LSUIn_valid ), .Z(\LSU/_0279_ ) );
BUF_X1 \LSU/_1610_ ( .A(_EXU_io_LSUIn_bits_wen ), .Z(\LSU/_0277_ ) );
BUF_X1 \LSU/_1611_ ( .A(_EXU_io_LSUIn_bits_ren ), .Z(\LSU/_0212_ ) );
BUF_X1 \LSU/_1612_ ( .A(\LSU/_0418_ ), .Z(_LSU_io_master_wlast ) );
BUF_X1 \LSU/_1613_ ( .A(\_LSU_io_master_awaddr [0] ), .Z(\LSU/_0316_ ) );
BUF_X1 \LSU/_1614_ ( .A(\_LSU_io_master_awaddr [1] ), .Z(\LSU/_0327_ ) );
BUF_X1 \LSU/_1615_ ( .A(\LSU/_0420_ ), .Z(\_LSU_io_master_wstrb [0] ) );
BUF_X1 \LSU/_1616_ ( .A(\LSU/_0004_ ), .Z(\LSU/_0009_ ) );
BUF_X1 \LSU/_1617_ ( .A(\LSU/_0003_ ), .Z(\LSU/_0008_ ) );
BUF_X1 \LSU/_1618_ ( .A(\LSU/_0421_ ), .Z(\_LSU_io_master_wstrb [1] ) );
BUF_X1 \LSU/_1619_ ( .A(\LSU/_0422_ ), .Z(\_LSU_io_master_wstrb [2] ) );
BUF_X1 \LSU/_1620_ ( .A(\LSU/_0423_ ), .Z(\_LSU_io_master_wstrb [3] ) );
BUF_X1 \LSU/_1621_ ( .A(\LSU/in_wdata [0] ), .Z(\LSU/_0145_ ) );
BUF_X1 \LSU/_1622_ ( .A(\LSU/_0386_ ), .Z(\_LSU_io_master_wdata [0] ) );
BUF_X1 \LSU/_1623_ ( .A(\LSU/in_wdata [1] ), .Z(\LSU/_0156_ ) );
BUF_X1 \LSU/_1624_ ( .A(\LSU/_0397_ ), .Z(\_LSU_io_master_wdata [1] ) );
BUF_X1 \LSU/_1625_ ( .A(\LSU/in_wdata [2] ), .Z(\LSU/_0167_ ) );
BUF_X1 \LSU/_1626_ ( .A(\LSU/_0408_ ), .Z(\_LSU_io_master_wdata [2] ) );
BUF_X1 \LSU/_1627_ ( .A(\LSU/in_wdata [3] ), .Z(\LSU/_0170_ ) );
BUF_X1 \LSU/_1628_ ( .A(\LSU/_0411_ ), .Z(\_LSU_io_master_wdata [3] ) );
BUF_X1 \LSU/_1629_ ( .A(\LSU/in_wdata [4] ), .Z(\LSU/_0171_ ) );
BUF_X1 \LSU/_1630_ ( .A(\LSU/_0412_ ), .Z(\_LSU_io_master_wdata [4] ) );
BUF_X1 \LSU/_1631_ ( .A(\LSU/in_wdata [5] ), .Z(\LSU/_0172_ ) );
BUF_X1 \LSU/_1632_ ( .A(\LSU/_0413_ ), .Z(\_LSU_io_master_wdata [5] ) );
BUF_X1 \LSU/_1633_ ( .A(\LSU/in_wdata [6] ), .Z(\LSU/_0173_ ) );
BUF_X1 \LSU/_1634_ ( .A(\LSU/_0414_ ), .Z(\_LSU_io_master_wdata [6] ) );
BUF_X1 \LSU/_1635_ ( .A(\LSU/in_wdata [7] ), .Z(\LSU/_0174_ ) );
BUF_X1 \LSU/_1636_ ( .A(\LSU/_0415_ ), .Z(\_LSU_io_master_wdata [7] ) );
BUF_X1 \LSU/_1637_ ( .A(\LSU/in_wdata [8] ), .Z(\LSU/_0175_ ) );
BUF_X1 \LSU/_1638_ ( .A(\LSU/_0416_ ), .Z(\_LSU_io_master_wdata [8] ) );
BUF_X1 \LSU/_1639_ ( .A(\LSU/in_wdata [9] ), .Z(\LSU/_0176_ ) );
BUF_X1 \LSU/_1640_ ( .A(\LSU/_0417_ ), .Z(\_LSU_io_master_wdata [9] ) );
BUF_X1 \LSU/_1641_ ( .A(\LSU/in_wdata [10] ), .Z(\LSU/_0146_ ) );
BUF_X1 \LSU/_1642_ ( .A(\LSU/_0387_ ), .Z(\_LSU_io_master_wdata [10] ) );
BUF_X1 \LSU/_1643_ ( .A(\LSU/in_wdata [11] ), .Z(\LSU/_0147_ ) );
BUF_X1 \LSU/_1644_ ( .A(\LSU/_0388_ ), .Z(\_LSU_io_master_wdata [11] ) );
BUF_X1 \LSU/_1645_ ( .A(\LSU/in_wdata [12] ), .Z(\LSU/_0148_ ) );
BUF_X1 \LSU/_1646_ ( .A(\LSU/_0389_ ), .Z(\_LSU_io_master_wdata [12] ) );
BUF_X1 \LSU/_1647_ ( .A(\LSU/in_wdata [13] ), .Z(\LSU/_0149_ ) );
BUF_X1 \LSU/_1648_ ( .A(\LSU/_0390_ ), .Z(\_LSU_io_master_wdata [13] ) );
BUF_X1 \LSU/_1649_ ( .A(\LSU/in_wdata [14] ), .Z(\LSU/_0150_ ) );
BUF_X1 \LSU/_1650_ ( .A(\LSU/_0391_ ), .Z(\_LSU_io_master_wdata [14] ) );
BUF_X1 \LSU/_1651_ ( .A(\LSU/in_wdata [15] ), .Z(\LSU/_0151_ ) );
BUF_X1 \LSU/_1652_ ( .A(\LSU/_0392_ ), .Z(\_LSU_io_master_wdata [15] ) );
BUF_X1 \LSU/_1653_ ( .A(\LSU/in_wdata [16] ), .Z(\LSU/_0152_ ) );
BUF_X1 \LSU/_1654_ ( .A(\LSU/_0393_ ), .Z(\_LSU_io_master_wdata [16] ) );
BUF_X1 \LSU/_1655_ ( .A(\LSU/in_wdata [17] ), .Z(\LSU/_0153_ ) );
BUF_X1 \LSU/_1656_ ( .A(\LSU/_0394_ ), .Z(\_LSU_io_master_wdata [17] ) );
BUF_X1 \LSU/_1657_ ( .A(\LSU/in_wdata [18] ), .Z(\LSU/_0154_ ) );
BUF_X1 \LSU/_1658_ ( .A(\LSU/_0395_ ), .Z(\_LSU_io_master_wdata [18] ) );
BUF_X1 \LSU/_1659_ ( .A(\LSU/in_wdata [19] ), .Z(\LSU/_0155_ ) );
BUF_X1 \LSU/_1660_ ( .A(\LSU/_0396_ ), .Z(\_LSU_io_master_wdata [19] ) );
BUF_X1 \LSU/_1661_ ( .A(\LSU/in_wdata [20] ), .Z(\LSU/_0157_ ) );
BUF_X1 \LSU/_1662_ ( .A(\LSU/_0398_ ), .Z(\_LSU_io_master_wdata [20] ) );
BUF_X1 \LSU/_1663_ ( .A(\LSU/in_wdata [21] ), .Z(\LSU/_0158_ ) );
BUF_X1 \LSU/_1664_ ( .A(\LSU/_0399_ ), .Z(\_LSU_io_master_wdata [21] ) );
BUF_X1 \LSU/_1665_ ( .A(\LSU/in_wdata [22] ), .Z(\LSU/_0159_ ) );
BUF_X1 \LSU/_1666_ ( .A(\LSU/_0400_ ), .Z(\_LSU_io_master_wdata [22] ) );
BUF_X1 \LSU/_1667_ ( .A(\LSU/in_wdata [23] ), .Z(\LSU/_0160_ ) );
BUF_X1 \LSU/_1668_ ( .A(\LSU/_0401_ ), .Z(\_LSU_io_master_wdata [23] ) );
BUF_X1 \LSU/_1669_ ( .A(\LSU/in_wdata [24] ), .Z(\LSU/_0161_ ) );
BUF_X1 \LSU/_1670_ ( .A(\LSU/_0402_ ), .Z(\_LSU_io_master_wdata [24] ) );
BUF_X1 \LSU/_1671_ ( .A(\LSU/in_wdata [25] ), .Z(\LSU/_0162_ ) );
BUF_X1 \LSU/_1672_ ( .A(\LSU/_0403_ ), .Z(\_LSU_io_master_wdata [25] ) );
BUF_X1 \LSU/_1673_ ( .A(\LSU/in_wdata [26] ), .Z(\LSU/_0163_ ) );
BUF_X1 \LSU/_1674_ ( .A(\LSU/_0404_ ), .Z(\_LSU_io_master_wdata [26] ) );
BUF_X1 \LSU/_1675_ ( .A(\LSU/in_wdata [27] ), .Z(\LSU/_0164_ ) );
BUF_X1 \LSU/_1676_ ( .A(\LSU/_0405_ ), .Z(\_LSU_io_master_wdata [27] ) );
BUF_X1 \LSU/_1677_ ( .A(\LSU/in_wdata [28] ), .Z(\LSU/_0165_ ) );
BUF_X1 \LSU/_1678_ ( .A(\LSU/_0406_ ), .Z(\_LSU_io_master_wdata [28] ) );
BUF_X1 \LSU/_1679_ ( .A(\LSU/in_wdata [29] ), .Z(\LSU/_0166_ ) );
BUF_X1 \LSU/_1680_ ( .A(\LSU/_0407_ ), .Z(\_LSU_io_master_wdata [29] ) );
BUF_X1 \LSU/_1681_ ( .A(\LSU/in_wdata [30] ), .Z(\LSU/_0168_ ) );
BUF_X1 \LSU/_1682_ ( .A(\LSU/_0409_ ), .Z(\_LSU_io_master_wdata [30] ) );
BUF_X1 \LSU/_1683_ ( .A(\LSU/in_wdata [31] ), .Z(\LSU/_0169_ ) );
BUF_X1 \LSU/_1684_ ( .A(\LSU/_0410_ ), .Z(\_LSU_io_master_wdata [31] ) );
BUF_X1 \LSU/_1685_ ( .A(\_AXI4Interconnect_io_fanIn_1_rdata [0] ), .Z(\LSU/_0352_ ) );
BUF_X1 \LSU/_1686_ ( .A(\_AXI4Interconnect_io_fanIn_1_rdata [1] ), .Z(\LSU/_0363_ ) );
BUF_X1 \LSU/_1687_ ( .A(\_AXI4Interconnect_io_fanIn_1_rdata [2] ), .Z(\LSU/_0374_ ) );
BUF_X1 \LSU/_1688_ ( .A(\_AXI4Interconnect_io_fanIn_1_rdata [3] ), .Z(\LSU/_0377_ ) );
BUF_X1 \LSU/_1689_ ( .A(\_AXI4Interconnect_io_fanIn_1_rdata [4] ), .Z(\LSU/_0378_ ) );
BUF_X1 \LSU/_1690_ ( .A(\_AXI4Interconnect_io_fanIn_1_rdata [5] ), .Z(\LSU/_0379_ ) );
BUF_X1 \LSU/_1691_ ( .A(\_AXI4Interconnect_io_fanIn_1_rdata [6] ), .Z(\LSU/_0380_ ) );
BUF_X1 \LSU/_1692_ ( .A(\_LSU_io_out_bits_rdata [0] ), .Z(\LSU/_0424_ ) );
BUF_X1 \LSU/_1693_ ( .A(\LSU/_0112_ ), .Z(\LSU/_0952_ ) );
BUF_X1 \LSU/_1694_ ( .A(\_LSU_io_out_bits_rdata [1] ), .Z(\LSU/_0435_ ) );
BUF_X1 \LSU/_1695_ ( .A(\LSU/_0113_ ), .Z(\LSU/_0953_ ) );
BUF_X1 \LSU/_1696_ ( .A(\_LSU_io_out_bits_rdata [2] ), .Z(\LSU/_0446_ ) );
BUF_X1 \LSU/_1697_ ( .A(\LSU/_0114_ ), .Z(\LSU/_0954_ ) );
BUF_X1 \LSU/_1698_ ( .A(\_LSU_io_out_bits_rdata [3] ), .Z(\LSU/_0449_ ) );
BUF_X1 \LSU/_1699_ ( .A(\LSU/_0115_ ), .Z(\LSU/_0955_ ) );
BUF_X1 \LSU/_1700_ ( .A(\_LSU_io_out_bits_rdata [4] ), .Z(\LSU/_0450_ ) );
BUF_X1 \LSU/_1701_ ( .A(\LSU/_0116_ ), .Z(\LSU/_0956_ ) );
BUF_X1 \LSU/_1702_ ( .A(\_LSU_io_out_bits_rdata [5] ), .Z(\LSU/_0451_ ) );
BUF_X1 \LSU/_1703_ ( .A(\LSU/_0117_ ), .Z(\LSU/_0957_ ) );
BUF_X1 \LSU/_1704_ ( .A(\_LSU_io_out_bits_rdata [6] ), .Z(\LSU/_0452_ ) );
BUF_X1 \LSU/_1705_ ( .A(\LSU/_0118_ ), .Z(\LSU/_0958_ ) );
BUF_X1 \LSU/_1706_ ( .A(\_LSU_io_out_bits_rdata [7] ), .Z(\LSU/_0453_ ) );
BUF_X1 \LSU/_1707_ ( .A(\LSU/_0119_ ), .Z(\LSU/_0959_ ) );
BUF_X1 \LSU/_1708_ ( .A(\_LSU_io_out_bits_rdata [8] ), .Z(\LSU/_0454_ ) );
BUF_X1 \LSU/_1709_ ( .A(\LSU/_0120_ ), .Z(\LSU/_0960_ ) );
BUF_X1 \LSU/_1710_ ( .A(\_LSU_io_out_bits_rdata [9] ), .Z(\LSU/_0455_ ) );
BUF_X1 \LSU/_1711_ ( .A(\LSU/_0121_ ), .Z(\LSU/_0961_ ) );
BUF_X1 \LSU/_1712_ ( .A(\_LSU_io_out_bits_rdata [10] ), .Z(\LSU/_0425_ ) );
BUF_X1 \LSU/_1713_ ( .A(\LSU/_0122_ ), .Z(\LSU/_0962_ ) );
BUF_X1 \LSU/_1714_ ( .A(\_LSU_io_out_bits_rdata [11] ), .Z(\LSU/_0426_ ) );
BUF_X1 \LSU/_1715_ ( .A(\LSU/_0123_ ), .Z(\LSU/_0963_ ) );
BUF_X1 \LSU/_1716_ ( .A(\_LSU_io_out_bits_rdata [12] ), .Z(\LSU/_0427_ ) );
BUF_X1 \LSU/_1717_ ( .A(\LSU/_0124_ ), .Z(\LSU/_0964_ ) );
BUF_X1 \LSU/_1718_ ( .A(\_LSU_io_out_bits_rdata [13] ), .Z(\LSU/_0428_ ) );
BUF_X1 \LSU/_1719_ ( .A(\LSU/_0125_ ), .Z(\LSU/_0965_ ) );
BUF_X1 \LSU/_1720_ ( .A(\_LSU_io_out_bits_rdata [14] ), .Z(\LSU/_0429_ ) );
BUF_X1 \LSU/_1721_ ( .A(\LSU/_0126_ ), .Z(\LSU/_0966_ ) );
BUF_X1 \LSU/_1722_ ( .A(\_LSU_io_out_bits_rdata [15] ), .Z(\LSU/_0430_ ) );
BUF_X1 \LSU/_1723_ ( .A(\LSU/_0127_ ), .Z(\LSU/_0967_ ) );
BUF_X1 \LSU/_1724_ ( .A(\_LSU_io_out_bits_rdata [16] ), .Z(\LSU/_0431_ ) );
BUF_X1 \LSU/_1725_ ( .A(\LSU/_0128_ ), .Z(\LSU/_0968_ ) );
BUF_X1 \LSU/_1726_ ( .A(\_LSU_io_out_bits_rdata [17] ), .Z(\LSU/_0432_ ) );
BUF_X1 \LSU/_1727_ ( .A(\LSU/_0129_ ), .Z(\LSU/_0969_ ) );
BUF_X1 \LSU/_1728_ ( .A(\_LSU_io_out_bits_rdata [18] ), .Z(\LSU/_0433_ ) );
BUF_X1 \LSU/_1729_ ( .A(\LSU/_0130_ ), .Z(\LSU/_0970_ ) );
BUF_X1 \LSU/_1730_ ( .A(\_LSU_io_out_bits_rdata [19] ), .Z(\LSU/_0434_ ) );
BUF_X1 \LSU/_1731_ ( .A(\LSU/_0131_ ), .Z(\LSU/_0971_ ) );
BUF_X1 \LSU/_1732_ ( .A(\_LSU_io_out_bits_rdata [20] ), .Z(\LSU/_0436_ ) );
BUF_X1 \LSU/_1733_ ( .A(\LSU/_0132_ ), .Z(\LSU/_0972_ ) );
BUF_X1 \LSU/_1734_ ( .A(\_LSU_io_out_bits_rdata [21] ), .Z(\LSU/_0437_ ) );
BUF_X1 \LSU/_1735_ ( .A(\LSU/_0133_ ), .Z(\LSU/_0973_ ) );
BUF_X1 \LSU/_1736_ ( .A(\_LSU_io_out_bits_rdata [22] ), .Z(\LSU/_0438_ ) );
BUF_X1 \LSU/_1737_ ( .A(\LSU/_0134_ ), .Z(\LSU/_0974_ ) );
BUF_X1 \LSU/_1738_ ( .A(\_LSU_io_out_bits_rdata [23] ), .Z(\LSU/_0439_ ) );
BUF_X1 \LSU/_1739_ ( .A(\LSU/_0135_ ), .Z(\LSU/_0975_ ) );
BUF_X1 \LSU/_1740_ ( .A(\_LSU_io_out_bits_rdata [24] ), .Z(\LSU/_0440_ ) );
BUF_X1 \LSU/_1741_ ( .A(\LSU/_0136_ ), .Z(\LSU/_0976_ ) );
BUF_X1 \LSU/_1742_ ( .A(\_LSU_io_out_bits_rdata [25] ), .Z(\LSU/_0441_ ) );
BUF_X1 \LSU/_1743_ ( .A(\LSU/_0137_ ), .Z(\LSU/_0977_ ) );
BUF_X1 \LSU/_1744_ ( .A(\_LSU_io_out_bits_rdata [26] ), .Z(\LSU/_0442_ ) );
BUF_X1 \LSU/_1745_ ( .A(\LSU/_0138_ ), .Z(\LSU/_0978_ ) );
BUF_X1 \LSU/_1746_ ( .A(\_LSU_io_out_bits_rdata [27] ), .Z(\LSU/_0443_ ) );
BUF_X1 \LSU/_1747_ ( .A(\LSU/_0139_ ), .Z(\LSU/_0979_ ) );
BUF_X1 \LSU/_1748_ ( .A(\_LSU_io_out_bits_rdata [28] ), .Z(\LSU/_0444_ ) );
BUF_X1 \LSU/_1749_ ( .A(\LSU/_0140_ ), .Z(\LSU/_0980_ ) );
BUF_X1 \LSU/_1750_ ( .A(\_LSU_io_out_bits_rdata [29] ), .Z(\LSU/_0445_ ) );
BUF_X1 \LSU/_1751_ ( .A(\LSU/_0141_ ), .Z(\LSU/_0981_ ) );
BUF_X1 \LSU/_1752_ ( .A(\_LSU_io_out_bits_rdata [30] ), .Z(\LSU/_0447_ ) );
BUF_X1 \LSU/_1753_ ( .A(\LSU/_0142_ ), .Z(\LSU/_0982_ ) );
BUF_X1 \LSU/_1754_ ( .A(\_LSU_io_out_bits_rdata [31] ), .Z(\LSU/_0448_ ) );
BUF_X1 \LSU/_1755_ ( .A(\LSU/_0143_ ), .Z(\LSU/_0983_ ) );
BUF_X1 \LSU/_1756_ ( .A(\_EXU_io_LSUIn_bits_memOp [0] ), .Z(\LSU/_0177_ ) );
BUF_X1 \LSU/_1757_ ( .A(\LSU/_0013_ ), .Z(\LSU/_0853_ ) );
BUF_X1 \LSU/_1758_ ( .A(\_EXU_io_LSUIn_bits_memOp [1] ), .Z(\LSU/_0178_ ) );
BUF_X1 \LSU/_1759_ ( .A(\LSU/_0014_ ), .Z(\LSU/_0854_ ) );
BUF_X1 \LSU/_1760_ ( .A(\_EXU_io_LSUIn_bits_memOp [2] ), .Z(\LSU/_0179_ ) );
BUF_X1 \LSU/_1761_ ( .A(\LSU/_0015_ ), .Z(\LSU/_0855_ ) );
BUF_X1 \LSU/_1762_ ( .A(\_EXU_io_LSUIn_bits_raddr [0] ), .Z(\LSU/_0180_ ) );
BUF_X1 \LSU/_1763_ ( .A(\LSU/_0016_ ), .Z(\LSU/_0856_ ) );
BUF_X1 \LSU/_1764_ ( .A(\_EXU_io_LSUIn_bits_raddr [1] ), .Z(\LSU/_0191_ ) );
BUF_X1 \LSU/_1765_ ( .A(\LSU/_0017_ ), .Z(\LSU/_0857_ ) );
BUF_X1 \LSU/_1766_ ( .A(\_EXU_io_LSUIn_bits_raddr [2] ), .Z(\LSU/_0202_ ) );
BUF_X1 \LSU/_1767_ ( .A(\_LSU_io_master_araddr [2] ), .Z(\LSU/_0302_ ) );
BUF_X1 \LSU/_1768_ ( .A(\LSU/_0018_ ), .Z(\LSU/_0858_ ) );
BUF_X1 \LSU/_1769_ ( .A(\_EXU_io_LSUIn_bits_raddr [3] ), .Z(\LSU/_0205_ ) );
BUF_X1 \LSU/_1770_ ( .A(\_LSU_io_master_araddr [3] ), .Z(\LSU/_0305_ ) );
BUF_X1 \LSU/_1771_ ( .A(\LSU/_0019_ ), .Z(\LSU/_0859_ ) );
BUF_X1 \LSU/_1772_ ( .A(\_EXU_io_LSUIn_bits_raddr [4] ), .Z(\LSU/_0206_ ) );
BUF_X1 \LSU/_1773_ ( .A(\_LSU_io_master_araddr [4] ), .Z(\LSU/_0306_ ) );
BUF_X1 \LSU/_1774_ ( .A(\LSU/_0020_ ), .Z(\LSU/_0860_ ) );
BUF_X1 \LSU/_1775_ ( .A(\_EXU_io_LSUIn_bits_raddr [5] ), .Z(\LSU/_0207_ ) );
BUF_X1 \LSU/_1776_ ( .A(\_LSU_io_master_araddr [5] ), .Z(\LSU/_0307_ ) );
BUF_X1 \LSU/_1777_ ( .A(\LSU/_0021_ ), .Z(\LSU/_0861_ ) );
BUF_X1 \LSU/_1778_ ( .A(\_EXU_io_LSUIn_bits_raddr [6] ), .Z(\LSU/_0208_ ) );
BUF_X1 \LSU/_1779_ ( .A(\_LSU_io_master_araddr [6] ), .Z(\LSU/_0308_ ) );
BUF_X1 \LSU/_1780_ ( .A(\LSU/_0022_ ), .Z(\LSU/_0862_ ) );
BUF_X1 \LSU/_1781_ ( .A(\_EXU_io_LSUIn_bits_raddr [7] ), .Z(\LSU/_0209_ ) );
BUF_X1 \LSU/_1782_ ( .A(\_LSU_io_master_araddr [7] ), .Z(\LSU/_0309_ ) );
BUF_X1 \LSU/_1783_ ( .A(\LSU/_0023_ ), .Z(\LSU/_0863_ ) );
BUF_X1 \LSU/_1784_ ( .A(\_EXU_io_LSUIn_bits_raddr [8] ), .Z(\LSU/_0210_ ) );
BUF_X1 \LSU/_1785_ ( .A(\_LSU_io_master_araddr [8] ), .Z(\LSU/_0310_ ) );
BUF_X1 \LSU/_1786_ ( .A(\LSU/_0024_ ), .Z(\LSU/_0864_ ) );
BUF_X1 \LSU/_1787_ ( .A(\_EXU_io_LSUIn_bits_raddr [9] ), .Z(\LSU/_0211_ ) );
BUF_X1 \LSU/_1788_ ( .A(\_LSU_io_master_araddr [9] ), .Z(\LSU/_0311_ ) );
BUF_X1 \LSU/_1789_ ( .A(\LSU/_0025_ ), .Z(\LSU/_0865_ ) );
BUF_X1 \LSU/_1790_ ( .A(\_EXU_io_LSUIn_bits_raddr [10] ), .Z(\LSU/_0181_ ) );
BUF_X1 \LSU/_1791_ ( .A(\_LSU_io_master_araddr [10] ), .Z(\LSU/_0281_ ) );
BUF_X1 \LSU/_1792_ ( .A(\LSU/_0026_ ), .Z(\LSU/_0866_ ) );
BUF_X1 \LSU/_1793_ ( .A(\_EXU_io_LSUIn_bits_raddr [11] ), .Z(\LSU/_0182_ ) );
BUF_X1 \LSU/_1794_ ( .A(\_LSU_io_master_araddr [11] ), .Z(\LSU/_0282_ ) );
BUF_X1 \LSU/_1795_ ( .A(\LSU/_0027_ ), .Z(\LSU/_0867_ ) );
BUF_X1 \LSU/_1796_ ( .A(\_EXU_io_LSUIn_bits_raddr [12] ), .Z(\LSU/_0183_ ) );
BUF_X1 \LSU/_1797_ ( .A(\_LSU_io_master_araddr [12] ), .Z(\LSU/_0283_ ) );
BUF_X1 \LSU/_1798_ ( .A(\LSU/_0028_ ), .Z(\LSU/_0868_ ) );
BUF_X1 \LSU/_1799_ ( .A(\_EXU_io_LSUIn_bits_raddr [13] ), .Z(\LSU/_0184_ ) );
BUF_X1 \LSU/_1800_ ( .A(\_LSU_io_master_araddr [13] ), .Z(\LSU/_0284_ ) );
BUF_X1 \LSU/_1801_ ( .A(\LSU/_0029_ ), .Z(\LSU/_0869_ ) );
BUF_X1 \LSU/_1802_ ( .A(\_EXU_io_LSUIn_bits_raddr [14] ), .Z(\LSU/_0185_ ) );
BUF_X1 \LSU/_1803_ ( .A(\_LSU_io_master_araddr [14] ), .Z(\LSU/_0285_ ) );
BUF_X1 \LSU/_1804_ ( .A(\LSU/_0030_ ), .Z(\LSU/_0870_ ) );
BUF_X1 \LSU/_1805_ ( .A(\_EXU_io_LSUIn_bits_raddr [15] ), .Z(\LSU/_0186_ ) );
BUF_X1 \LSU/_1806_ ( .A(\_LSU_io_master_araddr [15] ), .Z(\LSU/_0286_ ) );
BUF_X1 \LSU/_1807_ ( .A(\LSU/_0031_ ), .Z(\LSU/_0871_ ) );
BUF_X1 \LSU/_1808_ ( .A(\_EXU_io_LSUIn_bits_raddr [16] ), .Z(\LSU/_0187_ ) );
BUF_X1 \LSU/_1809_ ( .A(\_LSU_io_master_araddr [16] ), .Z(\LSU/_0287_ ) );
BUF_X1 \LSU/_1810_ ( .A(\LSU/_0032_ ), .Z(\LSU/_0872_ ) );
BUF_X1 \LSU/_1811_ ( .A(\_EXU_io_LSUIn_bits_raddr [17] ), .Z(\LSU/_0188_ ) );
BUF_X1 \LSU/_1812_ ( .A(\_LSU_io_master_araddr [17] ), .Z(\LSU/_0288_ ) );
BUF_X1 \LSU/_1813_ ( .A(\LSU/_0033_ ), .Z(\LSU/_0873_ ) );
BUF_X1 \LSU/_1814_ ( .A(\_EXU_io_LSUIn_bits_raddr [18] ), .Z(\LSU/_0189_ ) );
BUF_X1 \LSU/_1815_ ( .A(\_LSU_io_master_araddr [18] ), .Z(\LSU/_0289_ ) );
BUF_X1 \LSU/_1816_ ( .A(\LSU/_0034_ ), .Z(\LSU/_0874_ ) );
BUF_X1 \LSU/_1817_ ( .A(\_EXU_io_LSUIn_bits_raddr [19] ), .Z(\LSU/_0190_ ) );
BUF_X1 \LSU/_1818_ ( .A(\_LSU_io_master_araddr [19] ), .Z(\LSU/_0290_ ) );
BUF_X1 \LSU/_1819_ ( .A(\LSU/_0035_ ), .Z(\LSU/_0875_ ) );
BUF_X1 \LSU/_1820_ ( .A(\_EXU_io_LSUIn_bits_raddr [20] ), .Z(\LSU/_0192_ ) );
BUF_X1 \LSU/_1821_ ( .A(\_LSU_io_master_araddr [20] ), .Z(\LSU/_0292_ ) );
BUF_X1 \LSU/_1822_ ( .A(\LSU/_0036_ ), .Z(\LSU/_0876_ ) );
BUF_X1 \LSU/_1823_ ( .A(\_EXU_io_LSUIn_bits_raddr [21] ), .Z(\LSU/_0193_ ) );
BUF_X1 \LSU/_1824_ ( .A(\_LSU_io_master_araddr [21] ), .Z(\LSU/_0293_ ) );
BUF_X1 \LSU/_1825_ ( .A(\LSU/_0037_ ), .Z(\LSU/_0877_ ) );
BUF_X1 \LSU/_1826_ ( .A(\_EXU_io_LSUIn_bits_raddr [22] ), .Z(\LSU/_0194_ ) );
BUF_X1 \LSU/_1827_ ( .A(\_LSU_io_master_araddr [22] ), .Z(\LSU/_0294_ ) );
BUF_X1 \LSU/_1828_ ( .A(\LSU/_0038_ ), .Z(\LSU/_0878_ ) );
BUF_X1 \LSU/_1829_ ( .A(\_EXU_io_LSUIn_bits_raddr [23] ), .Z(\LSU/_0195_ ) );
BUF_X1 \LSU/_1830_ ( .A(\_LSU_io_master_araddr [23] ), .Z(\LSU/_0295_ ) );
BUF_X1 \LSU/_1831_ ( .A(\LSU/_0039_ ), .Z(\LSU/_0879_ ) );
BUF_X1 \LSU/_1832_ ( .A(\_EXU_io_LSUIn_bits_raddr [24] ), .Z(\LSU/_0196_ ) );
BUF_X1 \LSU/_1833_ ( .A(\_LSU_io_master_araddr [24] ), .Z(\LSU/_0296_ ) );
BUF_X1 \LSU/_1834_ ( .A(\LSU/_0040_ ), .Z(\LSU/_0880_ ) );
BUF_X1 \LSU/_1835_ ( .A(\_EXU_io_LSUIn_bits_raddr [25] ), .Z(\LSU/_0197_ ) );
BUF_X1 \LSU/_1836_ ( .A(\_LSU_io_master_araddr [25] ), .Z(\LSU/_0297_ ) );
BUF_X1 \LSU/_1837_ ( .A(\LSU/_0041_ ), .Z(\LSU/_0881_ ) );
BUF_X1 \LSU/_1838_ ( .A(\_EXU_io_LSUIn_bits_raddr [26] ), .Z(\LSU/_0198_ ) );
BUF_X1 \LSU/_1839_ ( .A(\_LSU_io_master_araddr [26] ), .Z(\LSU/_0298_ ) );
BUF_X1 \LSU/_1840_ ( .A(\LSU/_0042_ ), .Z(\LSU/_0882_ ) );
BUF_X1 \LSU/_1841_ ( .A(\_EXU_io_LSUIn_bits_raddr [27] ), .Z(\LSU/_0199_ ) );
BUF_X1 \LSU/_1842_ ( .A(\_LSU_io_master_araddr [27] ), .Z(\LSU/_0299_ ) );
BUF_X1 \LSU/_1843_ ( .A(\LSU/_0043_ ), .Z(\LSU/_0883_ ) );
BUF_X1 \LSU/_1844_ ( .A(\_EXU_io_LSUIn_bits_raddr [28] ), .Z(\LSU/_0200_ ) );
BUF_X1 \LSU/_1845_ ( .A(\_LSU_io_master_araddr [28] ), .Z(\LSU/_0300_ ) );
BUF_X1 \LSU/_1846_ ( .A(\LSU/_0044_ ), .Z(\LSU/_0884_ ) );
BUF_X1 \LSU/_1847_ ( .A(\_EXU_io_LSUIn_bits_raddr [29] ), .Z(\LSU/_0201_ ) );
BUF_X1 \LSU/_1848_ ( .A(\_LSU_io_master_araddr [29] ), .Z(\LSU/_0301_ ) );
BUF_X1 \LSU/_1849_ ( .A(\LSU/_0045_ ), .Z(\LSU/_0885_ ) );
BUF_X1 \LSU/_1850_ ( .A(\_EXU_io_LSUIn_bits_raddr [30] ), .Z(\LSU/_0203_ ) );
BUF_X1 \LSU/_1851_ ( .A(\_LSU_io_master_araddr [30] ), .Z(\LSU/_0303_ ) );
BUF_X1 \LSU/_1852_ ( .A(\LSU/_0046_ ), .Z(\LSU/_0886_ ) );
BUF_X1 \LSU/_1853_ ( .A(\_EXU_io_LSUIn_bits_raddr [31] ), .Z(\LSU/_0204_ ) );
BUF_X1 \LSU/_1854_ ( .A(\_LSU_io_master_araddr [31] ), .Z(\LSU/_0304_ ) );
BUF_X1 \LSU/_1855_ ( .A(\LSU/_0047_ ), .Z(\LSU/_0887_ ) );
BUF_X1 \LSU/_1856_ ( .A(\_EXU_io_LSUIn_bits_waddr [0] ), .Z(\LSU/_0213_ ) );
BUF_X1 \LSU/_1857_ ( .A(\LSU/_0048_ ), .Z(\LSU/_0888_ ) );
BUF_X1 \LSU/_1858_ ( .A(\_EXU_io_LSUIn_bits_waddr [1] ), .Z(\LSU/_0224_ ) );
BUF_X1 \LSU/_1859_ ( .A(\LSU/_0049_ ), .Z(\LSU/_0889_ ) );
BUF_X1 \LSU/_1860_ ( .A(\_EXU_io_LSUIn_bits_waddr [2] ), .Z(\LSU/_0235_ ) );
BUF_X1 \LSU/_1861_ ( .A(\_LSU_io_master_awaddr [2] ), .Z(\LSU/_0338_ ) );
BUF_X1 \LSU/_1862_ ( .A(\LSU/_0050_ ), .Z(\LSU/_0890_ ) );
BUF_X1 \LSU/_1863_ ( .A(\_EXU_io_LSUIn_bits_waddr [3] ), .Z(\LSU/_0238_ ) );
BUF_X1 \LSU/_1864_ ( .A(\_LSU_io_master_awaddr [3] ), .Z(\LSU/_0341_ ) );
BUF_X1 \LSU/_1865_ ( .A(\LSU/_0051_ ), .Z(\LSU/_0891_ ) );
BUF_X1 \LSU/_1866_ ( .A(\_EXU_io_LSUIn_bits_waddr [4] ), .Z(\LSU/_0239_ ) );
BUF_X1 \LSU/_1867_ ( .A(\_LSU_io_master_awaddr [4] ), .Z(\LSU/_0342_ ) );
BUF_X1 \LSU/_1868_ ( .A(\LSU/_0052_ ), .Z(\LSU/_0892_ ) );
BUF_X1 \LSU/_1869_ ( .A(\_EXU_io_LSUIn_bits_waddr [5] ), .Z(\LSU/_0240_ ) );
BUF_X1 \LSU/_1870_ ( .A(\_LSU_io_master_awaddr [5] ), .Z(\LSU/_0343_ ) );
BUF_X1 \LSU/_1871_ ( .A(\LSU/_0053_ ), .Z(\LSU/_0893_ ) );
BUF_X1 \LSU/_1872_ ( .A(\_EXU_io_LSUIn_bits_waddr [6] ), .Z(\LSU/_0241_ ) );
BUF_X1 \LSU/_1873_ ( .A(\_LSU_io_master_awaddr [6] ), .Z(\LSU/_0344_ ) );
BUF_X1 \LSU/_1874_ ( .A(\LSU/_0054_ ), .Z(\LSU/_0894_ ) );
BUF_X1 \LSU/_1875_ ( .A(\_EXU_io_LSUIn_bits_waddr [7] ), .Z(\LSU/_0242_ ) );
BUF_X1 \LSU/_1876_ ( .A(\_LSU_io_master_awaddr [7] ), .Z(\LSU/_0345_ ) );
BUF_X1 \LSU/_1877_ ( .A(\LSU/_0055_ ), .Z(\LSU/_0895_ ) );
BUF_X1 \LSU/_1878_ ( .A(\_EXU_io_LSUIn_bits_waddr [8] ), .Z(\LSU/_0243_ ) );
BUF_X1 \LSU/_1879_ ( .A(\_LSU_io_master_awaddr [8] ), .Z(\LSU/_0346_ ) );
BUF_X1 \LSU/_1880_ ( .A(\LSU/_0056_ ), .Z(\LSU/_0896_ ) );
BUF_X1 \LSU/_1881_ ( .A(\_EXU_io_LSUIn_bits_waddr [9] ), .Z(\LSU/_0244_ ) );
BUF_X1 \LSU/_1882_ ( .A(\_LSU_io_master_awaddr [9] ), .Z(\LSU/_0347_ ) );
BUF_X1 \LSU/_1883_ ( .A(\LSU/_0057_ ), .Z(\LSU/_0897_ ) );
BUF_X1 \LSU/_1884_ ( .A(\_EXU_io_LSUIn_bits_waddr [10] ), .Z(\LSU/_0214_ ) );
BUF_X1 \LSU/_1885_ ( .A(\_LSU_io_master_awaddr [10] ), .Z(\LSU/_0317_ ) );
BUF_X1 \LSU/_1886_ ( .A(\LSU/_0058_ ), .Z(\LSU/_0898_ ) );
BUF_X1 \LSU/_1887_ ( .A(\_EXU_io_LSUIn_bits_waddr [11] ), .Z(\LSU/_0215_ ) );
BUF_X1 \LSU/_1888_ ( .A(\_LSU_io_master_awaddr [11] ), .Z(\LSU/_0318_ ) );
BUF_X1 \LSU/_1889_ ( .A(\LSU/_0059_ ), .Z(\LSU/_0899_ ) );
BUF_X1 \LSU/_1890_ ( .A(\_EXU_io_LSUIn_bits_waddr [12] ), .Z(\LSU/_0216_ ) );
BUF_X1 \LSU/_1891_ ( .A(\_LSU_io_master_awaddr [12] ), .Z(\LSU/_0319_ ) );
BUF_X1 \LSU/_1892_ ( .A(\LSU/_0060_ ), .Z(\LSU/_0900_ ) );
BUF_X1 \LSU/_1893_ ( .A(\_EXU_io_LSUIn_bits_waddr [13] ), .Z(\LSU/_0217_ ) );
BUF_X1 \LSU/_1894_ ( .A(\_LSU_io_master_awaddr [13] ), .Z(\LSU/_0320_ ) );
BUF_X1 \LSU/_1895_ ( .A(\LSU/_0061_ ), .Z(\LSU/_0901_ ) );
BUF_X1 \LSU/_1896_ ( .A(\_EXU_io_LSUIn_bits_waddr [14] ), .Z(\LSU/_0218_ ) );
BUF_X1 \LSU/_1897_ ( .A(\_LSU_io_master_awaddr [14] ), .Z(\LSU/_0321_ ) );
BUF_X1 \LSU/_1898_ ( .A(\LSU/_0062_ ), .Z(\LSU/_0902_ ) );
BUF_X1 \LSU/_1899_ ( .A(\_EXU_io_LSUIn_bits_waddr [15] ), .Z(\LSU/_0219_ ) );
BUF_X1 \LSU/_1900_ ( .A(\_LSU_io_master_awaddr [15] ), .Z(\LSU/_0322_ ) );
BUF_X1 \LSU/_1901_ ( .A(\LSU/_0063_ ), .Z(\LSU/_0903_ ) );
BUF_X1 \LSU/_1902_ ( .A(\_EXU_io_LSUIn_bits_waddr [16] ), .Z(\LSU/_0220_ ) );
BUF_X1 \LSU/_1903_ ( .A(\_LSU_io_master_awaddr [16] ), .Z(\LSU/_0323_ ) );
BUF_X1 \LSU/_1904_ ( .A(\LSU/_0064_ ), .Z(\LSU/_0904_ ) );
BUF_X1 \LSU/_1905_ ( .A(\_EXU_io_LSUIn_bits_waddr [17] ), .Z(\LSU/_0221_ ) );
BUF_X1 \LSU/_1906_ ( .A(\_LSU_io_master_awaddr [17] ), .Z(\LSU/_0324_ ) );
BUF_X1 \LSU/_1907_ ( .A(\LSU/_0065_ ), .Z(\LSU/_0905_ ) );
BUF_X1 \LSU/_1908_ ( .A(\_EXU_io_LSUIn_bits_waddr [18] ), .Z(\LSU/_0222_ ) );
BUF_X1 \LSU/_1909_ ( .A(\_LSU_io_master_awaddr [18] ), .Z(\LSU/_0325_ ) );
BUF_X1 \LSU/_1910_ ( .A(\LSU/_0066_ ), .Z(\LSU/_0906_ ) );
BUF_X1 \LSU/_1911_ ( .A(\_EXU_io_LSUIn_bits_waddr [19] ), .Z(\LSU/_0223_ ) );
BUF_X1 \LSU/_1912_ ( .A(\_LSU_io_master_awaddr [19] ), .Z(\LSU/_0326_ ) );
BUF_X1 \LSU/_1913_ ( .A(\LSU/_0067_ ), .Z(\LSU/_0907_ ) );
BUF_X1 \LSU/_1914_ ( .A(\_EXU_io_LSUIn_bits_waddr [20] ), .Z(\LSU/_0225_ ) );
BUF_X1 \LSU/_1915_ ( .A(\_LSU_io_master_awaddr [20] ), .Z(\LSU/_0328_ ) );
BUF_X1 \LSU/_1916_ ( .A(\LSU/_0068_ ), .Z(\LSU/_0908_ ) );
BUF_X1 \LSU/_1917_ ( .A(\_EXU_io_LSUIn_bits_waddr [21] ), .Z(\LSU/_0226_ ) );
BUF_X1 \LSU/_1918_ ( .A(\_LSU_io_master_awaddr [21] ), .Z(\LSU/_0329_ ) );
BUF_X1 \LSU/_1919_ ( .A(\LSU/_0069_ ), .Z(\LSU/_0909_ ) );
BUF_X1 \LSU/_1920_ ( .A(\_EXU_io_LSUIn_bits_waddr [22] ), .Z(\LSU/_0227_ ) );
BUF_X1 \LSU/_1921_ ( .A(\_LSU_io_master_awaddr [22] ), .Z(\LSU/_0330_ ) );
BUF_X1 \LSU/_1922_ ( .A(\LSU/_0070_ ), .Z(\LSU/_0910_ ) );
BUF_X1 \LSU/_1923_ ( .A(\_EXU_io_LSUIn_bits_waddr [23] ), .Z(\LSU/_0228_ ) );
BUF_X1 \LSU/_1924_ ( .A(\_LSU_io_master_awaddr [23] ), .Z(\LSU/_0331_ ) );
BUF_X1 \LSU/_1925_ ( .A(\LSU/_0071_ ), .Z(\LSU/_0911_ ) );
BUF_X1 \LSU/_1926_ ( .A(\_EXU_io_LSUIn_bits_waddr [24] ), .Z(\LSU/_0229_ ) );
BUF_X1 \LSU/_1927_ ( .A(\_LSU_io_master_awaddr [24] ), .Z(\LSU/_0332_ ) );
BUF_X1 \LSU/_1928_ ( .A(\LSU/_0072_ ), .Z(\LSU/_0912_ ) );
BUF_X1 \LSU/_1929_ ( .A(\_EXU_io_LSUIn_bits_waddr [25] ), .Z(\LSU/_0230_ ) );
BUF_X1 \LSU/_1930_ ( .A(\_LSU_io_master_awaddr [25] ), .Z(\LSU/_0333_ ) );
BUF_X1 \LSU/_1931_ ( .A(\LSU/_0073_ ), .Z(\LSU/_0913_ ) );
BUF_X1 \LSU/_1932_ ( .A(\_EXU_io_LSUIn_bits_waddr [26] ), .Z(\LSU/_0231_ ) );
BUF_X1 \LSU/_1933_ ( .A(\_LSU_io_master_awaddr [26] ), .Z(\LSU/_0334_ ) );
BUF_X1 \LSU/_1934_ ( .A(\LSU/_0074_ ), .Z(\LSU/_0914_ ) );
BUF_X1 \LSU/_1935_ ( .A(\_EXU_io_LSUIn_bits_waddr [27] ), .Z(\LSU/_0232_ ) );
BUF_X1 \LSU/_1936_ ( .A(\_LSU_io_master_awaddr [27] ), .Z(\LSU/_0335_ ) );
BUF_X1 \LSU/_1937_ ( .A(\LSU/_0075_ ), .Z(\LSU/_0915_ ) );
BUF_X1 \LSU/_1938_ ( .A(\_EXU_io_LSUIn_bits_waddr [28] ), .Z(\LSU/_0233_ ) );
BUF_X1 \LSU/_1939_ ( .A(\_LSU_io_master_awaddr [28] ), .Z(\LSU/_0336_ ) );
BUF_X1 \LSU/_1940_ ( .A(\LSU/_0076_ ), .Z(\LSU/_0916_ ) );
BUF_X1 \LSU/_1941_ ( .A(\_EXU_io_LSUIn_bits_waddr [29] ), .Z(\LSU/_0234_ ) );
BUF_X1 \LSU/_1942_ ( .A(\_LSU_io_master_awaddr [29] ), .Z(\LSU/_0337_ ) );
BUF_X1 \LSU/_1943_ ( .A(\LSU/_0077_ ), .Z(\LSU/_0917_ ) );
BUF_X1 \LSU/_1944_ ( .A(\_EXU_io_LSUIn_bits_waddr [30] ), .Z(\LSU/_0236_ ) );
BUF_X1 \LSU/_1945_ ( .A(\_LSU_io_master_awaddr [30] ), .Z(\LSU/_0339_ ) );
BUF_X1 \LSU/_1946_ ( .A(\LSU/_0078_ ), .Z(\LSU/_0918_ ) );
BUF_X1 \LSU/_1947_ ( .A(\_EXU_io_LSUIn_bits_waddr [31] ), .Z(\LSU/_0237_ ) );
BUF_X1 \LSU/_1948_ ( .A(\_LSU_io_master_awaddr [31] ), .Z(\LSU/_0340_ ) );
BUF_X1 \LSU/_1949_ ( .A(\LSU/_0079_ ), .Z(\LSU/_0919_ ) );
BUF_X1 \LSU/_1950_ ( .A(\_EXU_io_LSUIn_bits_wdata [0] ), .Z(\LSU/_0245_ ) );
BUF_X1 \LSU/_1951_ ( .A(\LSU/_0080_ ), .Z(\LSU/_0920_ ) );
BUF_X1 \LSU/_1952_ ( .A(\_EXU_io_LSUIn_bits_wdata [1] ), .Z(\LSU/_0256_ ) );
BUF_X1 \LSU/_1953_ ( .A(\LSU/_0081_ ), .Z(\LSU/_0921_ ) );
BUF_X1 \LSU/_1954_ ( .A(\_EXU_io_LSUIn_bits_wdata [2] ), .Z(\LSU/_0267_ ) );
BUF_X1 \LSU/_1955_ ( .A(\LSU/_0082_ ), .Z(\LSU/_0922_ ) );
BUF_X1 \LSU/_1956_ ( .A(\_EXU_io_LSUIn_bits_wdata [3] ), .Z(\LSU/_0270_ ) );
BUF_X1 \LSU/_1957_ ( .A(\LSU/_0083_ ), .Z(\LSU/_0923_ ) );
BUF_X1 \LSU/_1958_ ( .A(\_EXU_io_LSUIn_bits_wdata [4] ), .Z(\LSU/_0271_ ) );
BUF_X1 \LSU/_1959_ ( .A(\LSU/_0084_ ), .Z(\LSU/_0924_ ) );
BUF_X1 \LSU/_1960_ ( .A(\_EXU_io_LSUIn_bits_wdata [5] ), .Z(\LSU/_0272_ ) );
BUF_X1 \LSU/_1961_ ( .A(\LSU/_0085_ ), .Z(\LSU/_0925_ ) );
BUF_X1 \LSU/_1962_ ( .A(\_EXU_io_LSUIn_bits_wdata [6] ), .Z(\LSU/_0273_ ) );
BUF_X1 \LSU/_1963_ ( .A(\LSU/_0086_ ), .Z(\LSU/_0926_ ) );
BUF_X1 \LSU/_1964_ ( .A(\_EXU_io_LSUIn_bits_wdata [7] ), .Z(\LSU/_0274_ ) );
BUF_X1 \LSU/_1965_ ( .A(\LSU/_0087_ ), .Z(\LSU/_0927_ ) );
BUF_X1 \LSU/_1966_ ( .A(\_EXU_io_LSUIn_bits_wdata [8] ), .Z(\LSU/_0275_ ) );
BUF_X1 \LSU/_1967_ ( .A(\LSU/_0088_ ), .Z(\LSU/_0928_ ) );
BUF_X1 \LSU/_1968_ ( .A(\_EXU_io_LSUIn_bits_wdata [9] ), .Z(\LSU/_0276_ ) );
BUF_X1 \LSU/_1969_ ( .A(\LSU/_0089_ ), .Z(\LSU/_0929_ ) );
BUF_X1 \LSU/_1970_ ( .A(\_EXU_io_LSUIn_bits_wdata [10] ), .Z(\LSU/_0246_ ) );
BUF_X1 \LSU/_1971_ ( .A(\LSU/_0090_ ), .Z(\LSU/_0930_ ) );
BUF_X1 \LSU/_1972_ ( .A(\_EXU_io_LSUIn_bits_wdata [11] ), .Z(\LSU/_0247_ ) );
BUF_X1 \LSU/_1973_ ( .A(\LSU/_0091_ ), .Z(\LSU/_0931_ ) );
BUF_X1 \LSU/_1974_ ( .A(\_EXU_io_LSUIn_bits_wdata [12] ), .Z(\LSU/_0248_ ) );
BUF_X1 \LSU/_1975_ ( .A(\LSU/_0092_ ), .Z(\LSU/_0932_ ) );
BUF_X1 \LSU/_1976_ ( .A(\_EXU_io_LSUIn_bits_wdata [13] ), .Z(\LSU/_0249_ ) );
BUF_X1 \LSU/_1977_ ( .A(\LSU/_0093_ ), .Z(\LSU/_0933_ ) );
BUF_X1 \LSU/_1978_ ( .A(\_EXU_io_LSUIn_bits_wdata [14] ), .Z(\LSU/_0250_ ) );
BUF_X1 \LSU/_1979_ ( .A(\LSU/_0094_ ), .Z(\LSU/_0934_ ) );
BUF_X1 \LSU/_1980_ ( .A(\_EXU_io_LSUIn_bits_wdata [15] ), .Z(\LSU/_0251_ ) );
BUF_X1 \LSU/_1981_ ( .A(\LSU/_0095_ ), .Z(\LSU/_0935_ ) );
BUF_X1 \LSU/_1982_ ( .A(\_EXU_io_LSUIn_bits_wdata [16] ), .Z(\LSU/_0252_ ) );
BUF_X1 \LSU/_1983_ ( .A(\LSU/_0096_ ), .Z(\LSU/_0936_ ) );
BUF_X1 \LSU/_1984_ ( .A(\_EXU_io_LSUIn_bits_wdata [17] ), .Z(\LSU/_0253_ ) );
BUF_X1 \LSU/_1985_ ( .A(\LSU/_0097_ ), .Z(\LSU/_0937_ ) );
BUF_X1 \LSU/_1986_ ( .A(\_EXU_io_LSUIn_bits_wdata [18] ), .Z(\LSU/_0254_ ) );
BUF_X1 \LSU/_1987_ ( .A(\LSU/_0098_ ), .Z(\LSU/_0938_ ) );
BUF_X1 \LSU/_1988_ ( .A(\_EXU_io_LSUIn_bits_wdata [19] ), .Z(\LSU/_0255_ ) );
BUF_X1 \LSU/_1989_ ( .A(\LSU/_0099_ ), .Z(\LSU/_0939_ ) );
BUF_X1 \LSU/_1990_ ( .A(\_EXU_io_LSUIn_bits_wdata [20] ), .Z(\LSU/_0257_ ) );
BUF_X1 \LSU/_1991_ ( .A(\LSU/_0100_ ), .Z(\LSU/_0940_ ) );
BUF_X1 \LSU/_1992_ ( .A(\_EXU_io_LSUIn_bits_wdata [21] ), .Z(\LSU/_0258_ ) );
BUF_X1 \LSU/_1993_ ( .A(\LSU/_0101_ ), .Z(\LSU/_0941_ ) );
BUF_X1 \LSU/_1994_ ( .A(\_EXU_io_LSUIn_bits_wdata [22] ), .Z(\LSU/_0259_ ) );
BUF_X1 \LSU/_1995_ ( .A(\LSU/_0102_ ), .Z(\LSU/_0942_ ) );
BUF_X1 \LSU/_1996_ ( .A(\_EXU_io_LSUIn_bits_wdata [23] ), .Z(\LSU/_0260_ ) );
BUF_X1 \LSU/_1997_ ( .A(\LSU/_0103_ ), .Z(\LSU/_0943_ ) );
BUF_X1 \LSU/_1998_ ( .A(\_EXU_io_LSUIn_bits_wdata [24] ), .Z(\LSU/_0261_ ) );
BUF_X1 \LSU/_1999_ ( .A(\LSU/_0104_ ), .Z(\LSU/_0944_ ) );
BUF_X1 \LSU/_2000_ ( .A(\_EXU_io_LSUIn_bits_wdata [25] ), .Z(\LSU/_0262_ ) );
BUF_X1 \LSU/_2001_ ( .A(\LSU/_0105_ ), .Z(\LSU/_0945_ ) );
BUF_X1 \LSU/_2002_ ( .A(\_EXU_io_LSUIn_bits_wdata [26] ), .Z(\LSU/_0263_ ) );
BUF_X1 \LSU/_2003_ ( .A(\LSU/_0106_ ), .Z(\LSU/_0946_ ) );
BUF_X1 \LSU/_2004_ ( .A(\_EXU_io_LSUIn_bits_wdata [27] ), .Z(\LSU/_0264_ ) );
BUF_X1 \LSU/_2005_ ( .A(\LSU/_0107_ ), .Z(\LSU/_0947_ ) );
BUF_X1 \LSU/_2006_ ( .A(\_EXU_io_LSUIn_bits_wdata [28] ), .Z(\LSU/_0265_ ) );
BUF_X1 \LSU/_2007_ ( .A(\LSU/_0108_ ), .Z(\LSU/_0948_ ) );
BUF_X1 \LSU/_2008_ ( .A(\_EXU_io_LSUIn_bits_wdata [29] ), .Z(\LSU/_0266_ ) );
BUF_X1 \LSU/_2009_ ( .A(\LSU/_0109_ ), .Z(\LSU/_0949_ ) );
BUF_X1 \LSU/_2010_ ( .A(\_EXU_io_LSUIn_bits_wdata [30] ), .Z(\LSU/_0268_ ) );
BUF_X1 \LSU/_2011_ ( .A(\LSU/_0110_ ), .Z(\LSU/_0950_ ) );
BUF_X1 \LSU/_2012_ ( .A(\_EXU_io_LSUIn_bits_wdata [31] ), .Z(\LSU/_0269_ ) );
BUF_X1 \LSU/_2013_ ( .A(\LSU/_0111_ ), .Z(\LSU/_0951_ ) );
BUF_X1 \LSU/_2014_ ( .A(reset ), .Z(\LSU/_0716_ ) );
BUF_X1 \LSU/_2015_ ( .A(\LSU/_0010_ ), .Z(\LSU/_0850_ ) );
BUF_X1 \LSU/_2016_ ( .A(\LSU/_0011_ ), .Z(\LSU/_0851_ ) );
BUF_X1 \LSU/_2017_ ( .A(\LSU/_0012_ ), .Z(\LSU/_0852_ ) );
INV_X1 \RegFile/_4754_ ( .A(\RegFile/_0642_ ), .ZN(\RegFile/_0749_ ) );
AND2_X1 \RegFile/_4755_ ( .A1(\RegFile/_0749_ ), .A2(\RegFile/_0643_ ), .ZN(\RegFile/_0750_ ) );
CLKBUF_X2 \RegFile/_4756_ ( .A(\RegFile/_0750_ ), .Z(\RegFile/_0751_ ) );
INV_X1 \RegFile/_4757_ ( .A(\RegFile/_0641_ ), .ZN(\RegFile/_0752_ ) );
AND2_X2 \RegFile/_4758_ ( .A1(\RegFile/_0752_ ), .A2(\RegFile/_0640_ ), .ZN(\RegFile/_0753_ ) );
AND3_X1 \RegFile/_4759_ ( .A1(\RegFile/_0751_ ), .A2(\RegFile/_0753_ ), .A3(\RegFile/_3762_ ), .ZN(\RegFile/_0754_ ) );
NOR2_X1 \RegFile/_4760_ ( .A1(\RegFile/_0752_ ), .A2(\RegFile/_0640_ ), .ZN(\RegFile/_0755_ ) );
AND2_X1 \RegFile/_4761_ ( .A1(\RegFile/_0750_ ), .A2(\RegFile/_0755_ ), .ZN(\RegFile/_0756_ ) );
NOR2_X1 \RegFile/_4762_ ( .A1(\RegFile/_0749_ ), .A2(\RegFile/_0643_ ), .ZN(\RegFile/_0757_ ) );
AND2_X1 \RegFile/_4763_ ( .A1(\RegFile/_0753_ ), .A2(\RegFile/_0757_ ), .ZN(\RegFile/_0758_ ) );
BUF_X4 \RegFile/_4764_ ( .A(\RegFile/_0758_ ), .Z(\RegFile/_0759_ ) );
AOI221_X4 \RegFile/_4765_ ( .A(\RegFile/_0754_ ), .B1(\RegFile/_0756_ ), .B2(\RegFile/_3314_ ), .C1(\RegFile/_3634_ ), .C2(\RegFile/_0759_ ), .ZN(\RegFile/_0760_ ) );
BUF_X4 \RegFile/_4766_ ( .A(\RegFile/_0753_ ), .Z(\RegFile/_0761_ ) );
BUF_X4 \RegFile/_4767_ ( .A(\RegFile/_0761_ ), .Z(\RegFile/_0762_ ) );
AND2_X1 \RegFile/_4768_ ( .A1(\RegFile/_0643_ ), .A2(\RegFile/_0642_ ), .ZN(\RegFile/_0763_ ) );
BUF_X4 \RegFile/_4769_ ( .A(\RegFile/_0763_ ), .Z(\RegFile/_0764_ ) );
BUF_X4 \RegFile/_4770_ ( .A(\RegFile/_0764_ ), .Z(\RegFile/_0765_ ) );
BUF_X4 \RegFile/_4771_ ( .A(\RegFile/_0765_ ), .Z(\RegFile/_0766_ ) );
NAND3_X1 \RegFile/_4772_ ( .A1(\RegFile/_0762_ ), .A2(\RegFile/_3410_ ), .A3(\RegFile/_0766_ ), .ZN(\RegFile/_0767_ ) );
NOR2_X1 \RegFile/_4773_ ( .A1(\RegFile/_0641_ ), .A2(\RegFile/_0640_ ), .ZN(\RegFile/_0768_ ) );
BUF_X4 \RegFile/_4774_ ( .A(\RegFile/_0768_ ), .Z(\RegFile/_0769_ ) );
BUF_X4 \RegFile/_4775_ ( .A(\RegFile/_0769_ ), .Z(\RegFile/_0770_ ) );
NAND3_X1 \RegFile/_4776_ ( .A1(\RegFile/_0766_ ), .A2(\RegFile/_0770_ ), .A3(\RegFile/_3378_ ), .ZN(\RegFile/_0771_ ) );
BUF_X2 \RegFile/_4777_ ( .A(\RegFile/_0750_ ), .Z(\RegFile/_0772_ ) );
AND2_X1 \RegFile/_4778_ ( .A1(\RegFile/_0641_ ), .A2(\RegFile/_0640_ ), .ZN(\RegFile/_0773_ ) );
BUF_X2 \RegFile/_4779_ ( .A(\RegFile/_0773_ ), .Z(\RegFile/_0774_ ) );
BUF_X2 \RegFile/_4780_ ( .A(\RegFile/_0774_ ), .Z(\RegFile/_0775_ ) );
AND3_X1 \RegFile/_4781_ ( .A1(\RegFile/_0772_ ), .A2(\RegFile/_3346_ ), .A3(\RegFile/_0775_ ), .ZN(\RegFile/_0776_ ) );
NOR2_X2 \RegFile/_4782_ ( .A1(\RegFile/_0643_ ), .A2(\RegFile/_0642_ ), .ZN(\RegFile/_0777_ ) );
AND2_X1 \RegFile/_4783_ ( .A1(\RegFile/_0773_ ), .A2(\RegFile/_0777_ ), .ZN(\RegFile/_0778_ ) );
BUF_X4 \RegFile/_4784_ ( .A(\RegFile/_0778_ ), .Z(\RegFile/_0779_ ) );
BUF_X4 \RegFile/_4785_ ( .A(\RegFile/_0779_ ), .Z(\RegFile/_0780_ ) );
AOI21_X1 \RegFile/_4786_ ( .A(\RegFile/_0776_ ), .B1(\RegFile/_3570_ ), .B2(\RegFile/_0780_ ), .ZN(\RegFile/_0781_ ) );
AND4_X1 \RegFile/_4787_ ( .A1(\RegFile/_0760_ ), .A2(\RegFile/_0767_ ), .A3(\RegFile/_0771_ ), .A4(\RegFile/_0781_ ), .ZN(\RegFile/_0782_ ) );
BUF_X4 \RegFile/_4788_ ( .A(\RegFile/_0755_ ), .Z(\RegFile/_0783_ ) );
BUF_X2 \RegFile/_4789_ ( .A(\RegFile/_0783_ ), .Z(\RegFile/_0784_ ) );
BUF_X4 \RegFile/_4790_ ( .A(\RegFile/_0784_ ), .Z(\RegFile/_0785_ ) );
BUF_X4 \RegFile/_4791_ ( .A(\RegFile/_0777_ ), .Z(\RegFile/_0786_ ) );
BUF_X4 \RegFile/_4792_ ( .A(\RegFile/_0786_ ), .Z(\RegFile/_0787_ ) );
NAND3_X1 \RegFile/_4793_ ( .A1(\RegFile/_0785_ ), .A2(\RegFile/_3538_ ), .A3(\RegFile/_0787_ ), .ZN(\RegFile/_0788_ ) );
AND2_X2 \RegFile/_4794_ ( .A1(\RegFile/_0755_ ), .A2(\RegFile/_0763_ ), .ZN(\RegFile/_0789_ ) );
INV_X2 \RegFile/_4795_ ( .A(\RegFile/_0789_ ), .ZN(\RegFile/_0790_ ) );
BUF_X2 \RegFile/_4796_ ( .A(\RegFile/_0790_ ), .Z(\RegFile/_0791_ ) );
OAI21_X1 \RegFile/_4797_ ( .A(\RegFile/_0788_ ), .B1(\RegFile/_0791_ ), .B2(\RegFile/_0111_ ), .ZN(\RegFile/_0792_ ) );
BUF_X2 \RegFile/_4798_ ( .A(\RegFile/_0772_ ), .Z(\RegFile/_0793_ ) );
BUF_X4 \RegFile/_4799_ ( .A(\RegFile/_0769_ ), .Z(\RegFile/_0794_ ) );
NAND3_X1 \RegFile/_4800_ ( .A1(\RegFile/_0793_ ), .A2(\RegFile/_3730_ ), .A3(\RegFile/_0794_ ), .ZN(\RegFile/_0795_ ) );
CLKBUF_X2 \RegFile/_4801_ ( .A(\RegFile/_0753_ ), .Z(\RegFile/_0796_ ) );
BUF_X4 \RegFile/_4802_ ( .A(\RegFile/_0777_ ), .Z(\RegFile/_0797_ ) );
NAND3_X1 \RegFile/_4803_ ( .A1(\RegFile/_0796_ ), .A2(\RegFile/_3506_ ), .A3(\RegFile/_0797_ ), .ZN(\RegFile/_0798_ ) );
BUF_X4 \RegFile/_4804_ ( .A(\RegFile/_0757_ ), .Z(\RegFile/_0799_ ) );
BUF_X4 \RegFile/_4805_ ( .A(\RegFile/_0799_ ), .Z(\RegFile/_0800_ ) );
BUF_X4 \RegFile/_4806_ ( .A(\RegFile/_0800_ ), .Z(\RegFile/_0801_ ) );
BUF_X4 \RegFile/_4807_ ( .A(\RegFile/_0768_ ), .Z(\RegFile/_0802_ ) );
NAND3_X1 \RegFile/_4808_ ( .A1(\RegFile/_0801_ ), .A2(\RegFile/_3602_ ), .A3(\RegFile/_0802_ ), .ZN(\RegFile/_0803_ ) );
NAND3_X1 \RegFile/_4809_ ( .A1(\RegFile/_0801_ ), .A2(\RegFile/_0784_ ), .A3(\RegFile/_3666_ ), .ZN(\RegFile/_0804_ ) );
NAND4_X1 \RegFile/_4810_ ( .A1(\RegFile/_0795_ ), .A2(\RegFile/_0798_ ), .A3(\RegFile/_0803_ ), .A4(\RegFile/_0804_ ), .ZN(\RegFile/_0805_ ) );
AND2_X1 \RegFile/_4811_ ( .A1(\RegFile/_0764_ ), .A2(\RegFile/_0774_ ), .ZN(\RegFile/_0806_ ) );
BUF_X4 \RegFile/_4812_ ( .A(\RegFile/_0806_ ), .Z(\RegFile/_0807_ ) );
BUF_X2 \RegFile/_4813_ ( .A(\RegFile/_0800_ ), .Z(\RegFile/_0808_ ) );
AND3_X1 \RegFile/_4814_ ( .A1(\RegFile/_0808_ ), .A2(\RegFile/_3698_ ), .A3(\RegFile/_0775_ ), .ZN(\RegFile/_0809_ ) );
NOR4_X1 \RegFile/_4815_ ( .A1(\RegFile/_0792_ ), .A2(\RegFile/_0805_ ), .A3(\RegFile/_0807_ ), .A4(\RegFile/_0809_ ), .ZN(\RegFile/_0810_ ) );
BUF_X4 \RegFile/_4816_ ( .A(\RegFile/_0807_ ), .Z(\RegFile/_0811_ ) );
BUF_X4 \RegFile/_4817_ ( .A(\RegFile/_0811_ ), .Z(\RegFile/_0812_ ) );
AOI22_X1 \RegFile/_4818_ ( .A1(\RegFile/_0782_ ), .A2(\RegFile/_0810_ ), .B1(\RegFile/_0110_ ), .B2(\RegFile/_0812_ ), .ZN(\RegFile/_0648_ ) );
INV_X1 \RegFile/_4819_ ( .A(\RegFile/_0806_ ), .ZN(\RegFile/_0813_ ) );
CLKBUF_X2 \RegFile/_4820_ ( .A(\RegFile/_0813_ ), .Z(\RegFile/_0814_ ) );
AND2_X1 \RegFile/_4821_ ( .A1(\RegFile/_0799_ ), .A2(\RegFile/_0755_ ), .ZN(\RegFile/_0815_ ) );
INV_X1 \RegFile/_4822_ ( .A(\RegFile/_0815_ ), .ZN(\RegFile/_0816_ ) );
INV_X1 \RegFile/_4823_ ( .A(\RegFile/_3677_ ), .ZN(\RegFile/_0817_ ) );
OAI22_X1 \RegFile/_4824_ ( .A1(\RegFile/_0816_ ), .A2(\RegFile/_0817_ ), .B1(\RegFile/_0790_ ), .B2(\RegFile/_0113_ ), .ZN(\RegFile/_0818_ ) );
AND2_X2 \RegFile/_4825_ ( .A1(\RegFile/_0755_ ), .A2(\RegFile/_0777_ ), .ZN(\RegFile/_0819_ ) );
BUF_X4 \RegFile/_4826_ ( .A(\RegFile/_0819_ ), .Z(\RegFile/_0820_ ) );
AND2_X2 \RegFile/_4827_ ( .A1(\RegFile/_0753_ ), .A2(\RegFile/_0777_ ), .ZN(\RegFile/_0821_ ) );
BUF_X4 \RegFile/_4828_ ( .A(\RegFile/_0821_ ), .Z(\RegFile/_0822_ ) );
AOI221_X4 \RegFile/_4829_ ( .A(\RegFile/_0818_ ), .B1(\RegFile/_3549_ ), .B2(\RegFile/_0820_ ), .C1(\RegFile/_3517_ ), .C2(\RegFile/_0822_ ), .ZN(\RegFile/_0823_ ) );
BUF_X4 \RegFile/_4830_ ( .A(\RegFile/_0772_ ), .Z(\RegFile/_0824_ ) );
BUF_X4 \RegFile/_4831_ ( .A(\RegFile/_0824_ ), .Z(\RegFile/_0825_ ) );
NAND3_X1 \RegFile/_4832_ ( .A1(\RegFile/_0825_ ), .A2(\RegFile/_3741_ ), .A3(\RegFile/_0770_ ), .ZN(\RegFile/_0826_ ) );
AND2_X2 \RegFile/_4833_ ( .A1(\RegFile/_0772_ ), .A2(\RegFile/_0753_ ), .ZN(\RegFile/_0827_ ) );
BUF_X4 \RegFile/_4834_ ( .A(\RegFile/_0827_ ), .Z(\RegFile/_0828_ ) );
BUF_X4 \RegFile/_4835_ ( .A(\RegFile/_0759_ ), .Z(\RegFile/_0829_ ) );
AOI22_X1 \RegFile/_4836_ ( .A1(\RegFile/_3773_ ), .A2(\RegFile/_0828_ ), .B1(\RegFile/_0829_ ), .B2(\RegFile/_3645_ ), .ZN(\RegFile/_0830_ ) );
AND4_X1 \RegFile/_4837_ ( .A1(\RegFile/_0814_ ), .A2(\RegFile/_0823_ ), .A3(\RegFile/_0826_ ), .A4(\RegFile/_0830_ ), .ZN(\RegFile/_0831_ ) );
BUF_X2 \RegFile/_4838_ ( .A(\RegFile/_0772_ ), .Z(\RegFile/_0832_ ) );
BUF_X4 \RegFile/_4839_ ( .A(\RegFile/_0832_ ), .Z(\RegFile/_0833_ ) );
BUF_X2 \RegFile/_4840_ ( .A(\RegFile/_0774_ ), .Z(\RegFile/_0834_ ) );
NAND3_X1 \RegFile/_4841_ ( .A1(\RegFile/_0833_ ), .A2(\RegFile/_3357_ ), .A3(\RegFile/_0834_ ), .ZN(\RegFile/_0835_ ) );
BUF_X4 \RegFile/_4842_ ( .A(\RegFile/_0769_ ), .Z(\RegFile/_0836_ ) );
NAND3_X1 \RegFile/_4843_ ( .A1(\RegFile/_0808_ ), .A2(\RegFile/_3613_ ), .A3(\RegFile/_0836_ ), .ZN(\RegFile/_0837_ ) );
INV_X1 \RegFile/_4844_ ( .A(\RegFile/_0780_ ), .ZN(\RegFile/_0838_ ) );
INV_X1 \RegFile/_4845_ ( .A(\RegFile/_3581_ ), .ZN(\RegFile/_0839_ ) );
OAI211_X2 \RegFile/_4846_ ( .A(\RegFile/_0835_ ), .B(\RegFile/_0837_ ), .C1(\RegFile/_0838_ ), .C2(\RegFile/_0839_ ), .ZN(\RegFile/_0840_ ) );
BUF_X2 \RegFile/_4847_ ( .A(\RegFile/_0753_ ), .Z(\RegFile/_0841_ ) );
BUF_X2 \RegFile/_4848_ ( .A(\RegFile/_0764_ ), .Z(\RegFile/_0842_ ) );
AND3_X1 \RegFile/_4849_ ( .A1(\RegFile/_0841_ ), .A2(\RegFile/_3421_ ), .A3(\RegFile/_0842_ ), .ZN(\RegFile/_0843_ ) );
CLKBUF_X2 \RegFile/_4850_ ( .A(\RegFile/_0772_ ), .Z(\RegFile/_0844_ ) );
AND3_X1 \RegFile/_4851_ ( .A1(\RegFile/_0844_ ), .A2(\RegFile/_0784_ ), .A3(\RegFile/_3325_ ), .ZN(\RegFile/_0845_ ) );
NAND3_X1 \RegFile/_4852_ ( .A1(\RegFile/_0765_ ), .A2(\RegFile/_0802_ ), .A3(\RegFile/_3389_ ), .ZN(\RegFile/_0846_ ) );
NAND2_X1 \RegFile/_4853_ ( .A1(\RegFile/_0800_ ), .A2(\RegFile/_0774_ ), .ZN(\RegFile/_0847_ ) );
BUF_X4 \RegFile/_4854_ ( .A(\RegFile/_0847_ ), .Z(\RegFile/_0848_ ) );
INV_X1 \RegFile/_4855_ ( .A(\RegFile/_3709_ ), .ZN(\RegFile/_0849_ ) );
OAI21_X1 \RegFile/_4856_ ( .A(\RegFile/_0846_ ), .B1(\RegFile/_0848_ ), .B2(\RegFile/_0849_ ), .ZN(\RegFile/_0850_ ) );
NOR4_X1 \RegFile/_4857_ ( .A1(\RegFile/_0840_ ), .A2(\RegFile/_0843_ ), .A3(\RegFile/_0845_ ), .A4(\RegFile/_0850_ ), .ZN(\RegFile/_0851_ ) );
AOI22_X1 \RegFile/_4858_ ( .A1(\RegFile/_0831_ ), .A2(\RegFile/_0851_ ), .B1(\RegFile/_0112_ ), .B2(\RegFile/_0812_ ), .ZN(\RegFile/_0659_ ) );
BUF_X4 \RegFile/_4859_ ( .A(\RegFile/_0765_ ), .Z(\RegFile/_0852_ ) );
NAND3_X1 \RegFile/_4860_ ( .A1(\RegFile/_0841_ ), .A2(\RegFile/_3432_ ), .A3(\RegFile/_0852_ ), .ZN(\RegFile/_0853_ ) );
NAND3_X1 \RegFile/_4861_ ( .A1(\RegFile/_0841_ ), .A2(\RegFile/_0808_ ), .A3(\RegFile/_3656_ ), .ZN(\RegFile/_0854_ ) );
BUF_X4 \RegFile/_4862_ ( .A(\RegFile/_0816_ ), .Z(\RegFile/_0855_ ) );
INV_X1 \RegFile/_4863_ ( .A(\RegFile/_3688_ ), .ZN(\RegFile/_0856_ ) );
OAI211_X2 \RegFile/_4864_ ( .A(\RegFile/_0853_ ), .B(\RegFile/_0854_ ), .C1(\RegFile/_0855_ ), .C2(\RegFile/_0856_ ), .ZN(\RegFile/_0857_ ) );
NAND3_X1 \RegFile/_4865_ ( .A1(\RegFile/_0833_ ), .A2(\RegFile/_3752_ ), .A3(\RegFile/_0836_ ), .ZN(\RegFile/_0858_ ) );
INV_X1 \RegFile/_4866_ ( .A(\RegFile/_3720_ ), .ZN(\RegFile/_0859_ ) );
OAI21_X1 \RegFile/_4867_ ( .A(\RegFile/_0858_ ), .B1(\RegFile/_0848_ ), .B2(\RegFile/_0859_ ), .ZN(\RegFile/_0860_ ) );
BUF_X2 \RegFile/_4868_ ( .A(\RegFile/_0753_ ), .Z(\RegFile/_0861_ ) );
AND3_X1 \RegFile/_4869_ ( .A1(\RegFile/_0793_ ), .A2(\RegFile/_0861_ ), .A3(\RegFile/_3784_ ), .ZN(\RegFile/_0862_ ) );
NOR4_X1 \RegFile/_4870_ ( .A1(\RegFile/_0857_ ), .A2(\RegFile/_0860_ ), .A3(\RegFile/_0807_ ), .A4(\RegFile/_0862_ ), .ZN(\RegFile/_0863_ ) );
CLKBUF_X2 \RegFile/_4871_ ( .A(\RegFile/_0772_ ), .Z(\RegFile/_0864_ ) );
AND3_X1 \RegFile/_4872_ ( .A1(\RegFile/_0864_ ), .A2(\RegFile/_3368_ ), .A3(\RegFile/_0775_ ), .ZN(\RegFile/_0865_ ) );
AOI21_X1 \RegFile/_4873_ ( .A(\RegFile/_0865_ ), .B1(\RegFile/_3336_ ), .B2(\RegFile/_0756_ ), .ZN(\RegFile/_0866_ ) );
INV_X1 \RegFile/_4874_ ( .A(\RegFile/_0115_ ), .ZN(\RegFile/_0867_ ) );
AND2_X1 \RegFile/_4875_ ( .A1(\RegFile/_0799_ ), .A2(\RegFile/_0768_ ), .ZN(\RegFile/_0868_ ) );
BUF_X4 \RegFile/_4876_ ( .A(\RegFile/_0868_ ), .Z(\RegFile/_0869_ ) );
BUF_X4 \RegFile/_4877_ ( .A(\RegFile/_0869_ ), .Z(\RegFile/_0870_ ) );
AOI22_X1 \RegFile/_4878_ ( .A1(\RegFile/_0867_ ), .A2(\RegFile/_0789_ ), .B1(\RegFile/_0870_ ), .B2(\RegFile/_3624_ ), .ZN(\RegFile/_0871_ ) );
AND2_X2 \RegFile/_4879_ ( .A1(\RegFile/_0764_ ), .A2(\RegFile/_0768_ ), .ZN(\RegFile/_0872_ ) );
AOI22_X1 \RegFile/_4880_ ( .A1(\RegFile/_0822_ ), .A2(\RegFile/_3528_ ), .B1(\RegFile/_0872_ ), .B2(\RegFile/_3400_ ), .ZN(\RegFile/_0873_ ) );
AOI22_X1 \RegFile/_4881_ ( .A1(\RegFile/_0820_ ), .A2(\RegFile/_3560_ ), .B1(\RegFile/_0780_ ), .B2(\RegFile/_3592_ ), .ZN(\RegFile/_0874_ ) );
AND4_X1 \RegFile/_4882_ ( .A1(\RegFile/_0866_ ), .A2(\RegFile/_0871_ ), .A3(\RegFile/_0873_ ), .A4(\RegFile/_0874_ ), .ZN(\RegFile/_0875_ ) );
AOI22_X1 \RegFile/_4883_ ( .A1(\RegFile/_0863_ ), .A2(\RegFile/_0875_ ), .B1(\RegFile/_0114_ ), .B2(\RegFile/_0812_ ), .ZN(\RegFile/_0670_ ) );
BUF_X2 \RegFile/_4884_ ( .A(\RegFile/_0755_ ), .Z(\RegFile/_0876_ ) );
NAND3_X1 \RegFile/_4885_ ( .A1(\RegFile/_0799_ ), .A2(\RegFile/_0876_ ), .A3(\RegFile/_3691_ ), .ZN(\RegFile/_0877_ ) );
OAI21_X1 \RegFile/_4886_ ( .A(\RegFile/_0877_ ), .B1(\RegFile/_0790_ ), .B2(\RegFile/_0117_ ), .ZN(\RegFile/_0878_ ) );
AOI221_X4 \RegFile/_4887_ ( .A(\RegFile/_0878_ ), .B1(\RegFile/_3563_ ), .B2(\RegFile/_0820_ ), .C1(\RegFile/_3531_ ), .C2(\RegFile/_0822_ ), .ZN(\RegFile/_0879_ ) );
NAND3_X1 \RegFile/_4888_ ( .A1(\RegFile/_0825_ ), .A2(\RegFile/_3755_ ), .A3(\RegFile/_0770_ ), .ZN(\RegFile/_0880_ ) );
AOI22_X1 \RegFile/_4889_ ( .A1(\RegFile/_3787_ ), .A2(\RegFile/_0828_ ), .B1(\RegFile/_0829_ ), .B2(\RegFile/_3659_ ), .ZN(\RegFile/_0881_ ) );
AND4_X1 \RegFile/_4890_ ( .A1(\RegFile/_0814_ ), .A2(\RegFile/_0879_ ), .A3(\RegFile/_0880_ ), .A4(\RegFile/_0881_ ), .ZN(\RegFile/_0882_ ) );
CLKBUF_X2 \RegFile/_4891_ ( .A(\RegFile/_0773_ ), .Z(\RegFile/_0883_ ) );
AND3_X1 \RegFile/_4892_ ( .A1(\RegFile/_0751_ ), .A2(\RegFile/_3371_ ), .A3(\RegFile/_0883_ ), .ZN(\RegFile/_0884_ ) );
AOI221_X4 \RegFile/_4893_ ( .A(\RegFile/_0884_ ), .B1(\RegFile/_3627_ ), .B2(\RegFile/_0869_ ), .C1(\RegFile/_3595_ ), .C2(\RegFile/_0780_ ), .ZN(\RegFile/_0885_ ) );
BUF_X2 \RegFile/_4894_ ( .A(\RegFile/_0783_ ), .Z(\RegFile/_0886_ ) );
AND3_X1 \RegFile/_4895_ ( .A1(\RegFile/_0832_ ), .A2(\RegFile/_0886_ ), .A3(\RegFile/_3339_ ), .ZN(\RegFile/_0887_ ) );
AND2_X2 \RegFile/_4896_ ( .A1(\RegFile/_0753_ ), .A2(\RegFile/_0764_ ), .ZN(\RegFile/_0888_ ) );
BUF_X4 \RegFile/_4897_ ( .A(\RegFile/_0888_ ), .Z(\RegFile/_0889_ ) );
AOI21_X1 \RegFile/_4898_ ( .A(\RegFile/_0887_ ), .B1(\RegFile/_3435_ ), .B2(\RegFile/_0889_ ), .ZN(\RegFile/_0890_ ) );
BUF_X4 \RegFile/_4899_ ( .A(\RegFile/_0769_ ), .Z(\RegFile/_0891_ ) );
NAND3_X1 \RegFile/_4900_ ( .A1(\RegFile/_0766_ ), .A2(\RegFile/_0891_ ), .A3(\RegFile/_3403_ ), .ZN(\RegFile/_0892_ ) );
BUF_X4 \RegFile/_4901_ ( .A(\RegFile/_0801_ ), .Z(\RegFile/_0893_ ) );
BUF_X2 \RegFile/_4902_ ( .A(\RegFile/_0774_ ), .Z(\RegFile/_0894_ ) );
NAND3_X1 \RegFile/_4903_ ( .A1(\RegFile/_0893_ ), .A2(\RegFile/_3723_ ), .A3(\RegFile/_0894_ ), .ZN(\RegFile/_0895_ ) );
AND4_X1 \RegFile/_4904_ ( .A1(\RegFile/_0885_ ), .A2(\RegFile/_0890_ ), .A3(\RegFile/_0892_ ), .A4(\RegFile/_0895_ ), .ZN(\RegFile/_0896_ ) );
AOI22_X1 \RegFile/_4905_ ( .A1(\RegFile/_0882_ ), .A2(\RegFile/_0896_ ), .B1(\RegFile/_0116_ ), .B2(\RegFile/_0812_ ), .ZN(\RegFile/_0673_ ) );
BUF_X4 \RegFile/_4906_ ( .A(\RegFile/_0801_ ), .Z(\RegFile/_0897_ ) );
BUF_X2 \RegFile/_4907_ ( .A(\RegFile/_0783_ ), .Z(\RegFile/_0898_ ) );
NAND3_X1 \RegFile/_4908_ ( .A1(\RegFile/_0897_ ), .A2(\RegFile/_0898_ ), .A3(\RegFile/_3692_ ), .ZN(\RegFile/_0899_ ) );
NAND3_X1 \RegFile/_4909_ ( .A1(\RegFile/_0841_ ), .A2(\RegFile/_3436_ ), .A3(\RegFile/_0852_ ), .ZN(\RegFile/_0900_ ) );
INV_X2 \RegFile/_4910_ ( .A(\RegFile/_0759_ ), .ZN(\RegFile/_0901_ ) );
INV_X1 \RegFile/_4911_ ( .A(\RegFile/_3660_ ), .ZN(\RegFile/_0902_ ) );
OAI211_X2 \RegFile/_4912_ ( .A(\RegFile/_0899_ ), .B(\RegFile/_0900_ ), .C1(\RegFile/_0901_ ), .C2(\RegFile/_0902_ ), .ZN(\RegFile/_0903_ ) );
NAND4_X1 \RegFile/_4913_ ( .A1(\RegFile/_0802_ ), .A2(\RegFile/_0643_ ), .A3(\RegFile/_0749_ ), .A4(\RegFile/_3756_ ), .ZN(\RegFile/_0904_ ) );
INV_X1 \RegFile/_4914_ ( .A(\RegFile/_3724_ ), .ZN(\RegFile/_0905_ ) );
OAI21_X1 \RegFile/_4915_ ( .A(\RegFile/_0904_ ), .B1(\RegFile/_0848_ ), .B2(\RegFile/_0905_ ), .ZN(\RegFile/_0906_ ) );
AND3_X1 \RegFile/_4916_ ( .A1(\RegFile/_0793_ ), .A2(\RegFile/_0861_ ), .A3(\RegFile/_3788_ ), .ZN(\RegFile/_0907_ ) );
NOR4_X1 \RegFile/_4917_ ( .A1(\RegFile/_0903_ ), .A2(\RegFile/_0811_ ), .A3(\RegFile/_0906_ ), .A4(\RegFile/_0907_ ), .ZN(\RegFile/_0908_ ) );
INV_X1 \RegFile/_4918_ ( .A(\RegFile/_0870_ ), .ZN(\RegFile/_0909_ ) );
INV_X1 \RegFile/_4919_ ( .A(\RegFile/_3628_ ), .ZN(\RegFile/_0910_ ) );
OAI22_X1 \RegFile/_4920_ ( .A1(\RegFile/_0791_ ), .A2(\RegFile/_0119_ ), .B1(\RegFile/_0909_ ), .B2(\RegFile/_0910_ ), .ZN(\RegFile/_0911_ ) );
BUF_X4 \RegFile/_4921_ ( .A(\RegFile/_0777_ ), .Z(\RegFile/_0912_ ) );
NAND3_X1 \RegFile/_4922_ ( .A1(\RegFile/_0834_ ), .A2(\RegFile/_0912_ ), .A3(\RegFile/_3596_ ), .ZN(\RegFile/_0913_ ) );
INV_X1 \RegFile/_4923_ ( .A(\RegFile/_0820_ ), .ZN(\RegFile/_0914_ ) );
INV_X1 \RegFile/_4924_ ( .A(\RegFile/_3564_ ), .ZN(\RegFile/_0915_ ) );
OAI21_X1 \RegFile/_4925_ ( .A(\RegFile/_0913_ ), .B1(\RegFile/_0914_ ), .B2(\RegFile/_0915_ ), .ZN(\RegFile/_0916_ ) );
NAND3_X1 \RegFile/_4926_ ( .A1(\RegFile/_0793_ ), .A2(\RegFile/_0898_ ), .A3(\RegFile/_3340_ ), .ZN(\RegFile/_0917_ ) );
BUF_X4 \RegFile/_4927_ ( .A(\RegFile/_0774_ ), .Z(\RegFile/_0918_ ) );
NAND3_X1 \RegFile/_4928_ ( .A1(\RegFile/_0793_ ), .A2(\RegFile/_3372_ ), .A3(\RegFile/_0918_ ), .ZN(\RegFile/_0919_ ) );
NAND2_X1 \RegFile/_4929_ ( .A1(\RegFile/_0917_ ), .A2(\RegFile/_0919_ ), .ZN(\RegFile/_0920_ ) );
NAND3_X1 \RegFile/_4930_ ( .A1(\RegFile/_0861_ ), .A2(\RegFile/_3532_ ), .A3(\RegFile/_0912_ ), .ZN(\RegFile/_0921_ ) );
NAND3_X1 \RegFile/_4931_ ( .A1(\RegFile/_0765_ ), .A2(\RegFile/_0794_ ), .A3(\RegFile/_3404_ ), .ZN(\RegFile/_0922_ ) );
NAND2_X1 \RegFile/_4932_ ( .A1(\RegFile/_0921_ ), .A2(\RegFile/_0922_ ), .ZN(\RegFile/_0923_ ) );
NOR4_X1 \RegFile/_4933_ ( .A1(\RegFile/_0911_ ), .A2(\RegFile/_0916_ ), .A3(\RegFile/_0920_ ), .A4(\RegFile/_0923_ ), .ZN(\RegFile/_0924_ ) );
AOI22_X1 \RegFile/_4934_ ( .A1(\RegFile/_0908_ ), .A2(\RegFile/_0924_ ), .B1(\RegFile/_0118_ ), .B2(\RegFile/_0812_ ), .ZN(\RegFile/_0674_ ) );
NAND3_X1 \RegFile/_4935_ ( .A1(\RegFile/_0799_ ), .A2(\RegFile/_0876_ ), .A3(\RegFile/_3693_ ), .ZN(\RegFile/_0925_ ) );
OAI21_X1 \RegFile/_4936_ ( .A(\RegFile/_0925_ ), .B1(\RegFile/_0790_ ), .B2(\RegFile/_0121_ ), .ZN(\RegFile/_0926_ ) );
AOI221_X4 \RegFile/_4937_ ( .A(\RegFile/_0926_ ), .B1(\RegFile/_3565_ ), .B2(\RegFile/_0820_ ), .C1(\RegFile/_3533_ ), .C2(\RegFile/_0822_ ), .ZN(\RegFile/_0927_ ) );
NAND3_X1 \RegFile/_4938_ ( .A1(\RegFile/_0825_ ), .A2(\RegFile/_3757_ ), .A3(\RegFile/_0770_ ), .ZN(\RegFile/_0928_ ) );
AOI22_X1 \RegFile/_4939_ ( .A1(\RegFile/_3789_ ), .A2(\RegFile/_0828_ ), .B1(\RegFile/_0829_ ), .B2(\RegFile/_3661_ ), .ZN(\RegFile/_0929_ ) );
AND4_X1 \RegFile/_4940_ ( .A1(\RegFile/_0814_ ), .A2(\RegFile/_0927_ ), .A3(\RegFile/_0928_ ), .A4(\RegFile/_0929_ ), .ZN(\RegFile/_0930_ ) );
AND3_X1 \RegFile/_4941_ ( .A1(\RegFile/_0751_ ), .A2(\RegFile/_3373_ ), .A3(\RegFile/_0883_ ), .ZN(\RegFile/_0931_ ) );
AOI221_X4 \RegFile/_4942_ ( .A(\RegFile/_0931_ ), .B1(\RegFile/_3629_ ), .B2(\RegFile/_0869_ ), .C1(\RegFile/_3597_ ), .C2(\RegFile/_0779_ ), .ZN(\RegFile/_0932_ ) );
AND3_X1 \RegFile/_4943_ ( .A1(\RegFile/_0832_ ), .A2(\RegFile/_0886_ ), .A3(\RegFile/_3341_ ), .ZN(\RegFile/_0933_ ) );
AOI21_X1 \RegFile/_4944_ ( .A(\RegFile/_0933_ ), .B1(\RegFile/_3437_ ), .B2(\RegFile/_0889_ ), .ZN(\RegFile/_0934_ ) );
NAND3_X1 \RegFile/_4945_ ( .A1(\RegFile/_0766_ ), .A2(\RegFile/_0891_ ), .A3(\RegFile/_3405_ ), .ZN(\RegFile/_0935_ ) );
NAND3_X1 \RegFile/_4946_ ( .A1(\RegFile/_0893_ ), .A2(\RegFile/_3725_ ), .A3(\RegFile/_0894_ ), .ZN(\RegFile/_0936_ ) );
AND4_X1 \RegFile/_4947_ ( .A1(\RegFile/_0932_ ), .A2(\RegFile/_0934_ ), .A3(\RegFile/_0935_ ), .A4(\RegFile/_0936_ ), .ZN(\RegFile/_0937_ ) );
AOI22_X1 \RegFile/_4948_ ( .A1(\RegFile/_0930_ ), .A2(\RegFile/_0937_ ), .B1(\RegFile/_0120_ ), .B2(\RegFile/_0812_ ), .ZN(\RegFile/_0675_ ) );
AND3_X1 \RegFile/_4949_ ( .A1(\RegFile/_0751_ ), .A2(\RegFile/_3374_ ), .A3(\RegFile/_0774_ ), .ZN(\RegFile/_0938_ ) );
AOI221_X4 \RegFile/_4950_ ( .A(\RegFile/_0938_ ), .B1(\RegFile/_3630_ ), .B2(\RegFile/_0869_ ), .C1(\RegFile/_3598_ ), .C2(\RegFile/_0780_ ), .ZN(\RegFile/_0939_ ) );
AND3_X1 \RegFile/_4951_ ( .A1(\RegFile/_0864_ ), .A2(\RegFile/_0784_ ), .A3(\RegFile/_3342_ ), .ZN(\RegFile/_0940_ ) );
AOI21_X1 \RegFile/_4952_ ( .A(\RegFile/_0940_ ), .B1(\RegFile/_3438_ ), .B2(\RegFile/_0889_ ), .ZN(\RegFile/_0941_ ) );
NAND3_X1 \RegFile/_4953_ ( .A1(\RegFile/_0766_ ), .A2(\RegFile/_0770_ ), .A3(\RegFile/_3406_ ), .ZN(\RegFile/_0942_ ) );
BUF_X4 \RegFile/_4954_ ( .A(\RegFile/_0775_ ), .Z(\RegFile/_0943_ ) );
NAND3_X1 \RegFile/_4955_ ( .A1(\RegFile/_0893_ ), .A2(\RegFile/_3726_ ), .A3(\RegFile/_0943_ ), .ZN(\RegFile/_0944_ ) );
AND4_X1 \RegFile/_4956_ ( .A1(\RegFile/_0939_ ), .A2(\RegFile/_0941_ ), .A3(\RegFile/_0942_ ), .A4(\RegFile/_0944_ ), .ZN(\RegFile/_0945_ ) );
AOI22_X1 \RegFile/_4957_ ( .A1(\RegFile/_3790_ ), .A2(\RegFile/_0828_ ), .B1(\RegFile/_0829_ ), .B2(\RegFile/_3662_ ), .ZN(\RegFile/_0946_ ) );
NAND3_X1 \RegFile/_4958_ ( .A1(\RegFile/_0761_ ), .A2(\RegFile/_3534_ ), .A3(\RegFile/_0786_ ), .ZN(\RegFile/_0947_ ) );
NAND3_X1 \RegFile/_4959_ ( .A1(\RegFile/_0801_ ), .A2(\RegFile/_0886_ ), .A3(\RegFile/_3694_ ), .ZN(\RegFile/_0948_ ) );
BUF_X2 \RegFile/_4960_ ( .A(\RegFile/_0783_ ), .Z(\RegFile/_0949_ ) );
NAND3_X1 \RegFile/_4961_ ( .A1(\RegFile/_0949_ ), .A2(\RegFile/_3566_ ), .A3(\RegFile/_0786_ ), .ZN(\RegFile/_0950_ ) );
INV_X1 \RegFile/_4962_ ( .A(\RegFile/_0123_ ), .ZN(\RegFile/_0951_ ) );
NAND3_X1 \RegFile/_4963_ ( .A1(\RegFile/_0783_ ), .A2(\RegFile/_0951_ ), .A3(\RegFile/_0765_ ), .ZN(\RegFile/_0952_ ) );
AND4_X1 \RegFile/_4964_ ( .A1(\RegFile/_0947_ ), .A2(\RegFile/_0948_ ), .A3(\RegFile/_0950_ ), .A4(\RegFile/_0952_ ), .ZN(\RegFile/_0953_ ) );
BUF_X4 \RegFile/_4965_ ( .A(\RegFile/_0824_ ), .Z(\RegFile/_0954_ ) );
BUF_X4 \RegFile/_4966_ ( .A(\RegFile/_0769_ ), .Z(\RegFile/_0955_ ) );
NAND3_X1 \RegFile/_4967_ ( .A1(\RegFile/_0954_ ), .A2(\RegFile/_3758_ ), .A3(\RegFile/_0955_ ), .ZN(\RegFile/_0956_ ) );
AND4_X1 \RegFile/_4968_ ( .A1(\RegFile/_0813_ ), .A2(\RegFile/_0946_ ), .A3(\RegFile/_0953_ ), .A4(\RegFile/_0956_ ), .ZN(\RegFile/_0957_ ) );
AOI22_X1 \RegFile/_4969_ ( .A1(\RegFile/_0945_ ), .A2(\RegFile/_0957_ ), .B1(\RegFile/_0122_ ), .B2(\RegFile/_0812_ ), .ZN(\RegFile/_0676_ ) );
AOI22_X1 \RegFile/_4970_ ( .A1(\RegFile/_3695_ ), .A2(\RegFile/_0815_ ), .B1(\RegFile/_0888_ ), .B2(\RegFile/_3439_ ), .ZN(\RegFile/_0958_ ) );
INV_X1 \RegFile/_4971_ ( .A(\RegFile/_3663_ ), .ZN(\RegFile/_0959_ ) );
OAI221_X1 \RegFile/_4972_ ( .A(\RegFile/_0958_ ), .B1(\RegFile/_0791_ ), .B2(\RegFile/_0125_ ), .C1(\RegFile/_0959_ ), .C2(\RegFile/_0901_ ), .ZN(\RegFile/_0960_ ) );
BUF_X2 \RegFile/_4973_ ( .A(\RegFile/_0772_ ), .Z(\RegFile/_0961_ ) );
AND3_X1 \RegFile/_4974_ ( .A1(\RegFile/_0961_ ), .A2(\RegFile/_3375_ ), .A3(\RegFile/_0894_ ), .ZN(\RegFile/_0962_ ) );
AND3_X1 \RegFile/_4975_ ( .A1(\RegFile/_0793_ ), .A2(\RegFile/_0898_ ), .A3(\RegFile/_3343_ ), .ZN(\RegFile/_0963_ ) );
NAND3_X1 \RegFile/_4976_ ( .A1(\RegFile/_0841_ ), .A2(\RegFile/_3535_ ), .A3(\RegFile/_0912_ ), .ZN(\RegFile/_0964_ ) );
NAND3_X1 \RegFile/_4977_ ( .A1(\RegFile/_0842_ ), .A2(\RegFile/_0794_ ), .A3(\RegFile/_3407_ ), .ZN(\RegFile/_0965_ ) );
NAND2_X1 \RegFile/_4978_ ( .A1(\RegFile/_0964_ ), .A2(\RegFile/_0965_ ), .ZN(\RegFile/_0966_ ) );
NOR4_X1 \RegFile/_4979_ ( .A1(\RegFile/_0960_ ), .A2(\RegFile/_0962_ ), .A3(\RegFile/_0963_ ), .A4(\RegFile/_0966_ ), .ZN(\RegFile/_0967_ ) );
AND3_X1 \RegFile/_4980_ ( .A1(\RegFile/_0876_ ), .A2(\RegFile/_3567_ ), .A3(\RegFile/_0777_ ), .ZN(\RegFile/_0968_ ) );
AOI221_X4 \RegFile/_4981_ ( .A(\RegFile/_0968_ ), .B1(\RegFile/_3599_ ), .B2(\RegFile/_0779_ ), .C1(\RegFile/_3631_ ), .C2(\RegFile/_0870_ ), .ZN(\RegFile/_0969_ ) );
NAND3_X1 \RegFile/_4982_ ( .A1(\RegFile/_0954_ ), .A2(\RegFile/_0762_ ), .A3(\RegFile/_3791_ ), .ZN(\RegFile/_0970_ ) );
AND3_X1 \RegFile/_4983_ ( .A1(\RegFile/_0800_ ), .A2(\RegFile/_3727_ ), .A3(\RegFile/_0774_ ), .ZN(\RegFile/_0971_ ) );
AND2_X1 \RegFile/_4984_ ( .A1(\RegFile/_0864_ ), .A2(\RegFile/_0769_ ), .ZN(\RegFile/_0972_ ) );
AOI21_X1 \RegFile/_4985_ ( .A(\RegFile/_0971_ ), .B1(\RegFile/_3759_ ), .B2(\RegFile/_0972_ ), .ZN(\RegFile/_0973_ ) );
AND4_X1 \RegFile/_4986_ ( .A1(\RegFile/_0813_ ), .A2(\RegFile/_0969_ ), .A3(\RegFile/_0970_ ), .A4(\RegFile/_0973_ ), .ZN(\RegFile/_0974_ ) );
AOI22_X1 \RegFile/_4987_ ( .A1(\RegFile/_0967_ ), .A2(\RegFile/_0974_ ), .B1(\RegFile/_0124_ ), .B2(\RegFile/_0812_ ), .ZN(\RegFile/_0677_ ) );
NAND3_X1 \RegFile/_4988_ ( .A1(\RegFile/_0762_ ), .A2(\RegFile/_3440_ ), .A3(\RegFile/_0852_ ), .ZN(\RegFile/_0975_ ) );
INV_X1 \RegFile/_4989_ ( .A(\RegFile/_3696_ ), .ZN(\RegFile/_0976_ ) );
INV_X1 \RegFile/_4990_ ( .A(\RegFile/_3664_ ), .ZN(\RegFile/_0977_ ) );
OAI221_X1 \RegFile/_4991_ ( .A(\RegFile/_0975_ ), .B1(\RegFile/_0855_ ), .B2(\RegFile/_0976_ ), .C1(\RegFile/_0977_ ), .C2(\RegFile/_0901_ ), .ZN(\RegFile/_0978_ ) );
NAND3_X1 \RegFile/_4992_ ( .A1(\RegFile/_0961_ ), .A2(\RegFile/_3760_ ), .A3(\RegFile/_0836_ ), .ZN(\RegFile/_0979_ ) );
NAND3_X1 \RegFile/_4993_ ( .A1(\RegFile/_0897_ ), .A2(\RegFile/_3728_ ), .A3(\RegFile/_0894_ ), .ZN(\RegFile/_0980_ ) );
NAND2_X1 \RegFile/_4994_ ( .A1(\RegFile/_0979_ ), .A2(\RegFile/_0980_ ), .ZN(\RegFile/_0981_ ) );
AND3_X1 \RegFile/_4995_ ( .A1(\RegFile/_0844_ ), .A2(\RegFile/_0861_ ), .A3(\RegFile/_3792_ ), .ZN(\RegFile/_0982_ ) );
NOR4_X1 \RegFile/_4996_ ( .A1(\RegFile/_0978_ ), .A2(\RegFile/_0981_ ), .A3(\RegFile/_0807_ ), .A4(\RegFile/_0982_ ), .ZN(\RegFile/_0983_ ) );
NAND3_X1 \RegFile/_4997_ ( .A1(\RegFile/_0897_ ), .A2(\RegFile/_3632_ ), .A3(\RegFile/_0955_ ), .ZN(\RegFile/_0984_ ) );
OAI21_X1 \RegFile/_4998_ ( .A(\RegFile/_0984_ ), .B1(\RegFile/_0791_ ), .B2(\RegFile/_0127_ ), .ZN(\RegFile/_0985_ ) );
NAND3_X1 \RegFile/_4999_ ( .A1(\RegFile/_0961_ ), .A2(\RegFile/_0785_ ), .A3(\RegFile/_3344_ ), .ZN(\RegFile/_0986_ ) );
NAND3_X1 \RegFile/_5000_ ( .A1(\RegFile/_0833_ ), .A2(\RegFile/_3376_ ), .A3(\RegFile/_0834_ ), .ZN(\RegFile/_0987_ ) );
NAND2_X1 \RegFile/_5001_ ( .A1(\RegFile/_0986_ ), .A2(\RegFile/_0987_ ), .ZN(\RegFile/_0988_ ) );
NAND3_X1 \RegFile/_5002_ ( .A1(\RegFile/_0861_ ), .A2(\RegFile/_3536_ ), .A3(\RegFile/_0912_ ), .ZN(\RegFile/_0989_ ) );
NAND3_X1 \RegFile/_5003_ ( .A1(\RegFile/_0842_ ), .A2(\RegFile/_0794_ ), .A3(\RegFile/_3408_ ), .ZN(\RegFile/_0990_ ) );
NAND2_X1 \RegFile/_5004_ ( .A1(\RegFile/_0989_ ), .A2(\RegFile/_0990_ ), .ZN(\RegFile/_0991_ ) );
NAND3_X1 \RegFile/_5005_ ( .A1(\RegFile/_0898_ ), .A2(\RegFile/_3568_ ), .A3(\RegFile/_0912_ ), .ZN(\RegFile/_0992_ ) );
NAND3_X1 \RegFile/_5006_ ( .A1(\RegFile/_0918_ ), .A2(\RegFile/_0797_ ), .A3(\RegFile/_3600_ ), .ZN(\RegFile/_0993_ ) );
NAND2_X1 \RegFile/_5007_ ( .A1(\RegFile/_0992_ ), .A2(\RegFile/_0993_ ), .ZN(\RegFile/_0994_ ) );
NOR4_X1 \RegFile/_5008_ ( .A1(\RegFile/_0985_ ), .A2(\RegFile/_0988_ ), .A3(\RegFile/_0991_ ), .A4(\RegFile/_0994_ ), .ZN(\RegFile/_0995_ ) );
AOI22_X1 \RegFile/_5009_ ( .A1(\RegFile/_0983_ ), .A2(\RegFile/_0995_ ), .B1(\RegFile/_0126_ ), .B2(\RegFile/_0812_ ), .ZN(\RegFile/_0678_ ) );
INV_X1 \RegFile/_5010_ ( .A(\RegFile/_3697_ ), .ZN(\RegFile/_0996_ ) );
OAI22_X1 \RegFile/_5011_ ( .A1(\RegFile/_0816_ ), .A2(\RegFile/_0996_ ), .B1(\RegFile/_0790_ ), .B2(\RegFile/_0065_ ), .ZN(\RegFile/_0997_ ) );
AOI221_X4 \RegFile/_5012_ ( .A(\RegFile/_0997_ ), .B1(\RegFile/_3569_ ), .B2(\RegFile/_0820_ ), .C1(\RegFile/_3537_ ), .C2(\RegFile/_0821_ ), .ZN(\RegFile/_0998_ ) );
NAND3_X1 \RegFile/_5013_ ( .A1(\RegFile/_0825_ ), .A2(\RegFile/_3761_ ), .A3(\RegFile/_0891_ ), .ZN(\RegFile/_0999_ ) );
AOI22_X1 \RegFile/_5014_ ( .A1(\RegFile/_3793_ ), .A2(\RegFile/_0828_ ), .B1(\RegFile/_0829_ ), .B2(\RegFile/_3665_ ), .ZN(\RegFile/_1000_ ) );
AND4_X1 \RegFile/_5015_ ( .A1(\RegFile/_0814_ ), .A2(\RegFile/_0998_ ), .A3(\RegFile/_0999_ ), .A4(\RegFile/_1000_ ), .ZN(\RegFile/_1001_ ) );
NAND3_X1 \RegFile/_5016_ ( .A1(\RegFile/_0833_ ), .A2(\RegFile/_3377_ ), .A3(\RegFile/_0918_ ), .ZN(\RegFile/_1002_ ) );
NAND3_X1 \RegFile/_5017_ ( .A1(\RegFile/_0834_ ), .A2(\RegFile/_0787_ ), .A3(\RegFile/_3601_ ), .ZN(\RegFile/_1003_ ) );
INV_X1 \RegFile/_5018_ ( .A(\RegFile/_3633_ ), .ZN(\RegFile/_1004_ ) );
OAI211_X2 \RegFile/_5019_ ( .A(\RegFile/_1002_ ), .B(\RegFile/_1003_ ), .C1(\RegFile/_0909_ ), .C2(\RegFile/_1004_ ), .ZN(\RegFile/_1005_ ) );
AND3_X1 \RegFile/_5020_ ( .A1(\RegFile/_0841_ ), .A2(\RegFile/_3441_ ), .A3(\RegFile/_0842_ ), .ZN(\RegFile/_1006_ ) );
AND3_X1 \RegFile/_5021_ ( .A1(\RegFile/_0844_ ), .A2(\RegFile/_0784_ ), .A3(\RegFile/_3345_ ), .ZN(\RegFile/_1007_ ) );
NAND3_X1 \RegFile/_5022_ ( .A1(\RegFile/_0765_ ), .A2(\RegFile/_0802_ ), .A3(\RegFile/_3409_ ), .ZN(\RegFile/_1008_ ) );
INV_X1 \RegFile/_5023_ ( .A(\RegFile/_3729_ ), .ZN(\RegFile/_1009_ ) );
OAI21_X1 \RegFile/_5024_ ( .A(\RegFile/_1008_ ), .B1(\RegFile/_0848_ ), .B2(\RegFile/_1009_ ), .ZN(\RegFile/_1010_ ) );
NOR4_X1 \RegFile/_5025_ ( .A1(\RegFile/_1005_ ), .A2(\RegFile/_1006_ ), .A3(\RegFile/_1007_ ), .A4(\RegFile/_1010_ ), .ZN(\RegFile/_1011_ ) );
AOI22_X1 \RegFile/_5026_ ( .A1(\RegFile/_1001_ ), .A2(\RegFile/_1011_ ), .B1(\RegFile/_0064_ ), .B2(\RegFile/_0812_ ), .ZN(\RegFile/_0679_ ) );
NAND3_X1 \RegFile/_5027_ ( .A1(\RegFile/_0762_ ), .A2(\RegFile/_3411_ ), .A3(\RegFile/_0852_ ), .ZN(\RegFile/_1012_ ) );
INV_X1 \RegFile/_5028_ ( .A(\RegFile/_3667_ ), .ZN(\RegFile/_1013_ ) );
INV_X1 \RegFile/_5029_ ( .A(\RegFile/_3635_ ), .ZN(\RegFile/_1014_ ) );
OAI221_X1 \RegFile/_5030_ ( .A(\RegFile/_1012_ ), .B1(\RegFile/_0855_ ), .B2(\RegFile/_1013_ ), .C1(\RegFile/_1014_ ), .C2(\RegFile/_0901_ ), .ZN(\RegFile/_1015_ ) );
NAND3_X1 \RegFile/_5031_ ( .A1(\RegFile/_0833_ ), .A2(\RegFile/_3731_ ), .A3(\RegFile/_0836_ ), .ZN(\RegFile/_1016_ ) );
NAND3_X1 \RegFile/_5032_ ( .A1(\RegFile/_0808_ ), .A2(\RegFile/_3699_ ), .A3(\RegFile/_0918_ ), .ZN(\RegFile/_1017_ ) );
NAND2_X1 \RegFile/_5033_ ( .A1(\RegFile/_1016_ ), .A2(\RegFile/_1017_ ), .ZN(\RegFile/_1018_ ) );
AND3_X1 \RegFile/_5034_ ( .A1(\RegFile/_0844_ ), .A2(\RegFile/_0796_ ), .A3(\RegFile/_3763_ ), .ZN(\RegFile/_1019_ ) );
NOR4_X1 \RegFile/_5035_ ( .A1(\RegFile/_1015_ ), .A2(\RegFile/_0811_ ), .A3(\RegFile/_1018_ ), .A4(\RegFile/_1019_ ), .ZN(\RegFile/_1020_ ) );
NAND3_X1 \RegFile/_5036_ ( .A1(\RegFile/_0897_ ), .A2(\RegFile/_3603_ ), .A3(\RegFile/_0836_ ), .ZN(\RegFile/_1021_ ) );
OAI21_X1 \RegFile/_5037_ ( .A(\RegFile/_1021_ ), .B1(\RegFile/_0791_ ), .B2(\RegFile/_0067_ ), .ZN(\RegFile/_1022_ ) );
NAND3_X1 \RegFile/_5038_ ( .A1(\RegFile/_0961_ ), .A2(\RegFile/_0785_ ), .A3(\RegFile/_3315_ ), .ZN(\RegFile/_1023_ ) );
NAND3_X1 \RegFile/_5039_ ( .A1(\RegFile/_0833_ ), .A2(\RegFile/_3347_ ), .A3(\RegFile/_0834_ ), .ZN(\RegFile/_1024_ ) );
NAND2_X1 \RegFile/_5040_ ( .A1(\RegFile/_1023_ ), .A2(\RegFile/_1024_ ), .ZN(\RegFile/_1025_ ) );
NAND3_X1 \RegFile/_5041_ ( .A1(\RegFile/_0861_ ), .A2(\RegFile/_3507_ ), .A3(\RegFile/_0912_ ), .ZN(\RegFile/_1026_ ) );
NAND3_X1 \RegFile/_5042_ ( .A1(\RegFile/_0842_ ), .A2(\RegFile/_0794_ ), .A3(\RegFile/_3379_ ), .ZN(\RegFile/_1027_ ) );
NAND2_X1 \RegFile/_5043_ ( .A1(\RegFile/_1026_ ), .A2(\RegFile/_1027_ ), .ZN(\RegFile/_1028_ ) );
NAND3_X1 \RegFile/_5044_ ( .A1(\RegFile/_0898_ ), .A2(\RegFile/_3539_ ), .A3(\RegFile/_0797_ ), .ZN(\RegFile/_1029_ ) );
NAND3_X1 \RegFile/_5045_ ( .A1(\RegFile/_0918_ ), .A2(\RegFile/_0797_ ), .A3(\RegFile/_3571_ ), .ZN(\RegFile/_1030_ ) );
NAND2_X1 \RegFile/_5046_ ( .A1(\RegFile/_1029_ ), .A2(\RegFile/_1030_ ), .ZN(\RegFile/_1031_ ) );
NOR4_X1 \RegFile/_5047_ ( .A1(\RegFile/_1022_ ), .A2(\RegFile/_1025_ ), .A3(\RegFile/_1028_ ), .A4(\RegFile/_1031_ ), .ZN(\RegFile/_1032_ ) );
BUF_X4 \RegFile/_5048_ ( .A(\RegFile/_0807_ ), .Z(\RegFile/_1033_ ) );
AOI22_X1 \RegFile/_5049_ ( .A1(\RegFile/_1020_ ), .A2(\RegFile/_1032_ ), .B1(\RegFile/_0066_ ), .B2(\RegFile/_1033_ ), .ZN(\RegFile/_0649_ ) );
NAND3_X1 \RegFile/_5050_ ( .A1(\RegFile/_0799_ ), .A2(\RegFile/_0876_ ), .A3(\RegFile/_3668_ ), .ZN(\RegFile/_1034_ ) );
OAI21_X1 \RegFile/_5051_ ( .A(\RegFile/_1034_ ), .B1(\RegFile/_0790_ ), .B2(\RegFile/_0069_ ), .ZN(\RegFile/_1035_ ) );
AOI221_X4 \RegFile/_5052_ ( .A(\RegFile/_1035_ ), .B1(\RegFile/_3540_ ), .B2(\RegFile/_0819_ ), .C1(\RegFile/_3508_ ), .C2(\RegFile/_0821_ ), .ZN(\RegFile/_1036_ ) );
NAND3_X1 \RegFile/_5053_ ( .A1(\RegFile/_0825_ ), .A2(\RegFile/_3732_ ), .A3(\RegFile/_0891_ ), .ZN(\RegFile/_1037_ ) );
AOI22_X1 \RegFile/_5054_ ( .A1(\RegFile/_3764_ ), .A2(\RegFile/_0827_ ), .B1(\RegFile/_0829_ ), .B2(\RegFile/_3636_ ), .ZN(\RegFile/_1038_ ) );
AND4_X1 \RegFile/_5055_ ( .A1(\RegFile/_0814_ ), .A2(\RegFile/_1036_ ), .A3(\RegFile/_1037_ ), .A4(\RegFile/_1038_ ), .ZN(\RegFile/_1039_ ) );
AND3_X1 \RegFile/_5056_ ( .A1(\RegFile/_0750_ ), .A2(\RegFile/_3348_ ), .A3(\RegFile/_0883_ ), .ZN(\RegFile/_1040_ ) );
AOI221_X4 \RegFile/_5057_ ( .A(\RegFile/_1040_ ), .B1(\RegFile/_3604_ ), .B2(\RegFile/_0869_ ), .C1(\RegFile/_3572_ ), .C2(\RegFile/_0779_ ), .ZN(\RegFile/_1041_ ) );
AND3_X1 \RegFile/_5058_ ( .A1(\RegFile/_0832_ ), .A2(\RegFile/_0886_ ), .A3(\RegFile/_3316_ ), .ZN(\RegFile/_1042_ ) );
AOI21_X1 \RegFile/_5059_ ( .A(\RegFile/_1042_ ), .B1(\RegFile/_3412_ ), .B2(\RegFile/_0889_ ), .ZN(\RegFile/_1043_ ) );
NAND3_X1 \RegFile/_5060_ ( .A1(\RegFile/_0766_ ), .A2(\RegFile/_0891_ ), .A3(\RegFile/_3380_ ), .ZN(\RegFile/_1044_ ) );
NAND3_X1 \RegFile/_5061_ ( .A1(\RegFile/_0897_ ), .A2(\RegFile/_3700_ ), .A3(\RegFile/_0894_ ), .ZN(\RegFile/_1045_ ) );
AND4_X1 \RegFile/_5062_ ( .A1(\RegFile/_1041_ ), .A2(\RegFile/_1043_ ), .A3(\RegFile/_1044_ ), .A4(\RegFile/_1045_ ), .ZN(\RegFile/_1046_ ) );
AOI22_X1 \RegFile/_5063_ ( .A1(\RegFile/_1039_ ), .A2(\RegFile/_1046_ ), .B1(\RegFile/_0068_ ), .B2(\RegFile/_1033_ ), .ZN(\RegFile/_0650_ ) );
NAND3_X1 \RegFile/_5064_ ( .A1(\RegFile/_0762_ ), .A2(\RegFile/_3413_ ), .A3(\RegFile/_0852_ ), .ZN(\RegFile/_1047_ ) );
INV_X1 \RegFile/_5065_ ( .A(\RegFile/_3669_ ), .ZN(\RegFile/_1048_ ) );
INV_X1 \RegFile/_5066_ ( .A(\RegFile/_3637_ ), .ZN(\RegFile/_1049_ ) );
OAI221_X1 \RegFile/_5067_ ( .A(\RegFile/_1047_ ), .B1(\RegFile/_0855_ ), .B2(\RegFile/_1048_ ), .C1(\RegFile/_1049_ ), .C2(\RegFile/_0901_ ), .ZN(\RegFile/_1050_ ) );
NAND4_X1 \RegFile/_5068_ ( .A1(\RegFile/_0802_ ), .A2(\RegFile/_0643_ ), .A3(\RegFile/_0749_ ), .A4(\RegFile/_3733_ ), .ZN(\RegFile/_1051_ ) );
INV_X1 \RegFile/_5069_ ( .A(\RegFile/_3701_ ), .ZN(\RegFile/_1052_ ) );
OAI21_X1 \RegFile/_5070_ ( .A(\RegFile/_1051_ ), .B1(\RegFile/_0848_ ), .B2(\RegFile/_1052_ ), .ZN(\RegFile/_1053_ ) );
AND3_X1 \RegFile/_5071_ ( .A1(\RegFile/_0844_ ), .A2(\RegFile/_0796_ ), .A3(\RegFile/_3765_ ), .ZN(\RegFile/_1054_ ) );
NOR4_X1 \RegFile/_5072_ ( .A1(\RegFile/_1050_ ), .A2(\RegFile/_0811_ ), .A3(\RegFile/_1053_ ), .A4(\RegFile/_1054_ ), .ZN(\RegFile/_1055_ ) );
INV_X1 \RegFile/_5073_ ( .A(\RegFile/_3605_ ), .ZN(\RegFile/_1056_ ) );
OAI22_X1 \RegFile/_5074_ ( .A1(\RegFile/_0791_ ), .A2(\RegFile/_0071_ ), .B1(\RegFile/_0909_ ), .B2(\RegFile/_1056_ ), .ZN(\RegFile/_1057_ ) );
NAND3_X1 \RegFile/_5075_ ( .A1(\RegFile/_0834_ ), .A2(\RegFile/_0912_ ), .A3(\RegFile/_3573_ ), .ZN(\RegFile/_1058_ ) );
INV_X1 \RegFile/_5076_ ( .A(\RegFile/_3541_ ), .ZN(\RegFile/_1059_ ) );
OAI21_X1 \RegFile/_5077_ ( .A(\RegFile/_1058_ ), .B1(\RegFile/_0914_ ), .B2(\RegFile/_1059_ ), .ZN(\RegFile/_1060_ ) );
NAND3_X1 \RegFile/_5078_ ( .A1(\RegFile/_0793_ ), .A2(\RegFile/_0898_ ), .A3(\RegFile/_3317_ ), .ZN(\RegFile/_1061_ ) );
NAND3_X1 \RegFile/_5079_ ( .A1(\RegFile/_0793_ ), .A2(\RegFile/_3349_ ), .A3(\RegFile/_0918_ ), .ZN(\RegFile/_1062_ ) );
NAND2_X1 \RegFile/_5080_ ( .A1(\RegFile/_1061_ ), .A2(\RegFile/_1062_ ), .ZN(\RegFile/_1063_ ) );
NAND3_X1 \RegFile/_5081_ ( .A1(\RegFile/_0861_ ), .A2(\RegFile/_3509_ ), .A3(\RegFile/_0797_ ), .ZN(\RegFile/_1064_ ) );
NAND3_X1 \RegFile/_5082_ ( .A1(\RegFile/_0765_ ), .A2(\RegFile/_0802_ ), .A3(\RegFile/_3381_ ), .ZN(\RegFile/_1065_ ) );
NAND2_X1 \RegFile/_5083_ ( .A1(\RegFile/_1064_ ), .A2(\RegFile/_1065_ ), .ZN(\RegFile/_1066_ ) );
NOR4_X1 \RegFile/_5084_ ( .A1(\RegFile/_1057_ ), .A2(\RegFile/_1060_ ), .A3(\RegFile/_1063_ ), .A4(\RegFile/_1066_ ), .ZN(\RegFile/_1067_ ) );
AOI22_X1 \RegFile/_5085_ ( .A1(\RegFile/_1055_ ), .A2(\RegFile/_1067_ ), .B1(\RegFile/_0070_ ), .B2(\RegFile/_1033_ ), .ZN(\RegFile/_0651_ ) );
NAND3_X1 \RegFile/_5086_ ( .A1(\RegFile/_0799_ ), .A2(\RegFile/_0876_ ), .A3(\RegFile/_3670_ ), .ZN(\RegFile/_1068_ ) );
OAI21_X1 \RegFile/_5087_ ( .A(\RegFile/_1068_ ), .B1(\RegFile/_0790_ ), .B2(\RegFile/_0073_ ), .ZN(\RegFile/_1069_ ) );
AOI221_X4 \RegFile/_5088_ ( .A(\RegFile/_1069_ ), .B1(\RegFile/_3542_ ), .B2(\RegFile/_0819_ ), .C1(\RegFile/_3510_ ), .C2(\RegFile/_0821_ ), .ZN(\RegFile/_1070_ ) );
NAND3_X1 \RegFile/_5089_ ( .A1(\RegFile/_0825_ ), .A2(\RegFile/_3734_ ), .A3(\RegFile/_0891_ ), .ZN(\RegFile/_1071_ ) );
AOI22_X1 \RegFile/_5090_ ( .A1(\RegFile/_3766_ ), .A2(\RegFile/_0827_ ), .B1(\RegFile/_0759_ ), .B2(\RegFile/_3638_ ), .ZN(\RegFile/_1072_ ) );
AND4_X1 \RegFile/_5091_ ( .A1(\RegFile/_0814_ ), .A2(\RegFile/_1070_ ), .A3(\RegFile/_1071_ ), .A4(\RegFile/_1072_ ), .ZN(\RegFile/_1073_ ) );
AND3_X1 \RegFile/_5092_ ( .A1(\RegFile/_0750_ ), .A2(\RegFile/_3350_ ), .A3(\RegFile/_0883_ ), .ZN(\RegFile/_1074_ ) );
AOI221_X4 \RegFile/_5093_ ( .A(\RegFile/_1074_ ), .B1(\RegFile/_3606_ ), .B2(\RegFile/_0869_ ), .C1(\RegFile/_3574_ ), .C2(\RegFile/_0779_ ), .ZN(\RegFile/_1075_ ) );
AND3_X1 \RegFile/_5094_ ( .A1(\RegFile/_0832_ ), .A2(\RegFile/_0886_ ), .A3(\RegFile/_3318_ ), .ZN(\RegFile/_1076_ ) );
AOI21_X1 \RegFile/_5095_ ( .A(\RegFile/_1076_ ), .B1(\RegFile/_3414_ ), .B2(\RegFile/_0889_ ), .ZN(\RegFile/_1077_ ) );
NAND3_X1 \RegFile/_5096_ ( .A1(\RegFile/_0852_ ), .A2(\RegFile/_0955_ ), .A3(\RegFile/_3382_ ), .ZN(\RegFile/_1078_ ) );
NAND3_X1 \RegFile/_5097_ ( .A1(\RegFile/_0897_ ), .A2(\RegFile/_3702_ ), .A3(\RegFile/_0894_ ), .ZN(\RegFile/_1079_ ) );
AND4_X1 \RegFile/_5098_ ( .A1(\RegFile/_1075_ ), .A2(\RegFile/_1077_ ), .A3(\RegFile/_1078_ ), .A4(\RegFile/_1079_ ), .ZN(\RegFile/_1080_ ) );
AOI22_X1 \RegFile/_5099_ ( .A1(\RegFile/_1073_ ), .A2(\RegFile/_1080_ ), .B1(\RegFile/_0072_ ), .B2(\RegFile/_1033_ ), .ZN(\RegFile/_0652_ ) );
NAND3_X1 \RegFile/_5100_ ( .A1(\RegFile/_0799_ ), .A2(\RegFile/_0876_ ), .A3(\RegFile/_3671_ ), .ZN(\RegFile/_1081_ ) );
OAI21_X1 \RegFile/_5101_ ( .A(\RegFile/_1081_ ), .B1(\RegFile/_0790_ ), .B2(\RegFile/_0075_ ), .ZN(\RegFile/_1082_ ) );
AOI221_X4 \RegFile/_5102_ ( .A(\RegFile/_1082_ ), .B1(\RegFile/_3543_ ), .B2(\RegFile/_0819_ ), .C1(\RegFile/_3511_ ), .C2(\RegFile/_0821_ ), .ZN(\RegFile/_1083_ ) );
NAND3_X1 \RegFile/_5103_ ( .A1(\RegFile/_0954_ ), .A2(\RegFile/_3735_ ), .A3(\RegFile/_0891_ ), .ZN(\RegFile/_1084_ ) );
AOI22_X1 \RegFile/_5104_ ( .A1(\RegFile/_3767_ ), .A2(\RegFile/_0827_ ), .B1(\RegFile/_0759_ ), .B2(\RegFile/_3639_ ), .ZN(\RegFile/_1085_ ) );
AND4_X1 \RegFile/_5105_ ( .A1(\RegFile/_0814_ ), .A2(\RegFile/_1083_ ), .A3(\RegFile/_1084_ ), .A4(\RegFile/_1085_ ), .ZN(\RegFile/_1086_ ) );
AND3_X1 \RegFile/_5106_ ( .A1(\RegFile/_0750_ ), .A2(\RegFile/_3351_ ), .A3(\RegFile/_0883_ ), .ZN(\RegFile/_1087_ ) );
AOI221_X4 \RegFile/_5107_ ( .A(\RegFile/_1087_ ), .B1(\RegFile/_3575_ ), .B2(\RegFile/_0779_ ), .C1(\RegFile/_3607_ ), .C2(\RegFile/_0870_ ), .ZN(\RegFile/_1088_ ) );
AND3_X1 \RegFile/_5108_ ( .A1(\RegFile/_0772_ ), .A2(\RegFile/_0886_ ), .A3(\RegFile/_3319_ ), .ZN(\RegFile/_1089_ ) );
AOI21_X1 \RegFile/_5109_ ( .A(\RegFile/_1089_ ), .B1(\RegFile/_3415_ ), .B2(\RegFile/_0889_ ), .ZN(\RegFile/_1090_ ) );
NAND3_X1 \RegFile/_5110_ ( .A1(\RegFile/_0852_ ), .A2(\RegFile/_0955_ ), .A3(\RegFile/_3383_ ), .ZN(\RegFile/_1091_ ) );
NAND3_X1 \RegFile/_5111_ ( .A1(\RegFile/_0897_ ), .A2(\RegFile/_3703_ ), .A3(\RegFile/_0894_ ), .ZN(\RegFile/_1092_ ) );
AND4_X1 \RegFile/_5112_ ( .A1(\RegFile/_1088_ ), .A2(\RegFile/_1090_ ), .A3(\RegFile/_1091_ ), .A4(\RegFile/_1092_ ), .ZN(\RegFile/_1093_ ) );
AOI22_X1 \RegFile/_5113_ ( .A1(\RegFile/_1086_ ), .A2(\RegFile/_1093_ ), .B1(\RegFile/_0074_ ), .B2(\RegFile/_1033_ ), .ZN(\RegFile/_0653_ ) );
NAND3_X1 \RegFile/_5114_ ( .A1(\RegFile/_0825_ ), .A2(\RegFile/_3352_ ), .A3(\RegFile/_0943_ ), .ZN(\RegFile/_1094_ ) );
NAND3_X1 \RegFile/_5115_ ( .A1(\RegFile/_0799_ ), .A2(\RegFile/_0876_ ), .A3(\RegFile/_3672_ ), .ZN(\RegFile/_1095_ ) );
INV_X1 \RegFile/_5116_ ( .A(\RegFile/_0888_ ), .ZN(\RegFile/_1096_ ) );
INV_X1 \RegFile/_5117_ ( .A(\RegFile/_3416_ ), .ZN(\RegFile/_1097_ ) );
OAI21_X1 \RegFile/_5118_ ( .A(\RegFile/_1095_ ), .B1(\RegFile/_1096_ ), .B2(\RegFile/_1097_ ), .ZN(\RegFile/_1098_ ) );
INV_X1 \RegFile/_5119_ ( .A(\RegFile/_0077_ ), .ZN(\RegFile/_1099_ ) );
AOI221_X4 \RegFile/_5120_ ( .A(\RegFile/_1098_ ), .B1(\RegFile/_1099_ ), .B2(\RegFile/_0789_ ), .C1(\RegFile/_3640_ ), .C2(\RegFile/_0759_ ), .ZN(\RegFile/_1100_ ) );
NAND3_X1 \RegFile/_5121_ ( .A1(\RegFile/_0954_ ), .A2(\RegFile/_0785_ ), .A3(\RegFile/_3320_ ), .ZN(\RegFile/_1101_ ) );
AOI22_X1 \RegFile/_5122_ ( .A1(\RegFile/_0822_ ), .A2(\RegFile/_3512_ ), .B1(\RegFile/_0872_ ), .B2(\RegFile/_3384_ ), .ZN(\RegFile/_1102_ ) );
AND4_X1 \RegFile/_5123_ ( .A1(\RegFile/_1094_ ), .A2(\RegFile/_1100_ ), .A3(\RegFile/_1101_ ), .A4(\RegFile/_1102_ ), .ZN(\RegFile/_1103_ ) );
NAND3_X1 \RegFile/_5124_ ( .A1(\RegFile/_0785_ ), .A2(\RegFile/_3544_ ), .A3(\RegFile/_0787_ ), .ZN(\RegFile/_1104_ ) );
NAND3_X1 \RegFile/_5125_ ( .A1(\RegFile/_0832_ ), .A2(\RegFile/_3736_ ), .A3(\RegFile/_0769_ ), .ZN(\RegFile/_1105_ ) );
NAND3_X1 \RegFile/_5126_ ( .A1(\RegFile/_0832_ ), .A2(\RegFile/_0761_ ), .A3(\RegFile/_3768_ ), .ZN(\RegFile/_1106_ ) );
NAND3_X1 \RegFile/_5127_ ( .A1(\RegFile/_0800_ ), .A2(\RegFile/_3704_ ), .A3(\RegFile/_0774_ ), .ZN(\RegFile/_1107_ ) );
AND4_X1 \RegFile/_5128_ ( .A1(\RegFile/_0813_ ), .A2(\RegFile/_1105_ ), .A3(\RegFile/_1106_ ), .A4(\RegFile/_1107_ ), .ZN(\RegFile/_1108_ ) );
NAND3_X1 \RegFile/_5129_ ( .A1(\RegFile/_0893_ ), .A2(\RegFile/_3608_ ), .A3(\RegFile/_0955_ ), .ZN(\RegFile/_1109_ ) );
NAND3_X1 \RegFile/_5130_ ( .A1(\RegFile/_0943_ ), .A2(\RegFile/_0787_ ), .A3(\RegFile/_3576_ ), .ZN(\RegFile/_1110_ ) );
AND4_X1 \RegFile/_5131_ ( .A1(\RegFile/_1104_ ), .A2(\RegFile/_1108_ ), .A3(\RegFile/_1109_ ), .A4(\RegFile/_1110_ ), .ZN(\RegFile/_1111_ ) );
AOI22_X1 \RegFile/_5132_ ( .A1(\RegFile/_1103_ ), .A2(\RegFile/_1111_ ), .B1(\RegFile/_0076_ ), .B2(\RegFile/_1033_ ), .ZN(\RegFile/_0654_ ) );
AND3_X1 \RegFile/_5133_ ( .A1(\RegFile/_0800_ ), .A2(\RegFile/_0876_ ), .A3(\RegFile/_3673_ ), .ZN(\RegFile/_1112_ ) );
AOI221_X4 \RegFile/_5134_ ( .A(\RegFile/_1112_ ), .B1(\RegFile/_0888_ ), .B2(\RegFile/_3417_ ), .C1(\RegFile/_3641_ ), .C2(\RegFile/_0759_ ), .ZN(\RegFile/_1113_ ) );
NAND3_X1 \RegFile/_5135_ ( .A1(\RegFile/_0954_ ), .A2(\RegFile/_0762_ ), .A3(\RegFile/_3769_ ), .ZN(\RegFile/_1114_ ) );
NAND3_X1 \RegFile/_5136_ ( .A1(\RegFile/_0824_ ), .A2(\RegFile/_3737_ ), .A3(\RegFile/_0769_ ), .ZN(\RegFile/_1115_ ) );
NAND3_X1 \RegFile/_5137_ ( .A1(\RegFile/_0801_ ), .A2(\RegFile/_3705_ ), .A3(\RegFile/_0775_ ), .ZN(\RegFile/_1116_ ) );
AND2_X1 \RegFile/_5138_ ( .A1(\RegFile/_1115_ ), .A2(\RegFile/_1116_ ), .ZN(\RegFile/_1117_ ) );
AND4_X1 \RegFile/_5139_ ( .A1(\RegFile/_0814_ ), .A2(\RegFile/_1113_ ), .A3(\RegFile/_1114_ ), .A4(\RegFile/_1117_ ), .ZN(\RegFile/_1118_ ) );
AND3_X1 \RegFile/_5140_ ( .A1(\RegFile/_0864_ ), .A2(\RegFile/_3353_ ), .A3(\RegFile/_0775_ ), .ZN(\RegFile/_1119_ ) );
AOI21_X1 \RegFile/_5141_ ( .A(\RegFile/_1119_ ), .B1(\RegFile/_3321_ ), .B2(\RegFile/_0756_ ), .ZN(\RegFile/_1120_ ) );
INV_X1 \RegFile/_5142_ ( .A(\RegFile/_0079_ ), .ZN(\RegFile/_1121_ ) );
AOI22_X1 \RegFile/_5143_ ( .A1(\RegFile/_1121_ ), .A2(\RegFile/_0789_ ), .B1(\RegFile/_0870_ ), .B2(\RegFile/_3609_ ), .ZN(\RegFile/_1122_ ) );
AOI22_X1 \RegFile/_5144_ ( .A1(\RegFile/_0822_ ), .A2(\RegFile/_3513_ ), .B1(\RegFile/_0872_ ), .B2(\RegFile/_3385_ ), .ZN(\RegFile/_1123_ ) );
AOI22_X1 \RegFile/_5145_ ( .A1(\RegFile/_0820_ ), .A2(\RegFile/_3545_ ), .B1(\RegFile/_0780_ ), .B2(\RegFile/_3577_ ), .ZN(\RegFile/_1124_ ) );
AND4_X1 \RegFile/_5146_ ( .A1(\RegFile/_1120_ ), .A2(\RegFile/_1122_ ), .A3(\RegFile/_1123_ ), .A4(\RegFile/_1124_ ), .ZN(\RegFile/_1125_ ) );
AOI22_X1 \RegFile/_5147_ ( .A1(\RegFile/_1118_ ), .A2(\RegFile/_1125_ ), .B1(\RegFile/_0078_ ), .B2(\RegFile/_1033_ ), .ZN(\RegFile/_0655_ ) );
NAND3_X1 \RegFile/_5148_ ( .A1(\RegFile/_0761_ ), .A2(\RegFile/_3514_ ), .A3(\RegFile/_0797_ ), .ZN(\RegFile/_1126_ ) );
OR2_X1 \RegFile/_5149_ ( .A1(\RegFile/_0791_ ), .A2(\RegFile/_0081_ ), .ZN(\RegFile/_1127_ ) );
NAND3_X1 \RegFile/_5150_ ( .A1(\RegFile/_0784_ ), .A2(\RegFile/_3546_ ), .A3(\RegFile/_0786_ ), .ZN(\RegFile/_1128_ ) );
NAND3_X1 \RegFile/_5151_ ( .A1(\RegFile/_0801_ ), .A2(\RegFile/_0949_ ), .A3(\RegFile/_3674_ ), .ZN(\RegFile/_1129_ ) );
AND4_X1 \RegFile/_5152_ ( .A1(\RegFile/_1126_ ), .A2(\RegFile/_1127_ ), .A3(\RegFile/_1128_ ), .A4(\RegFile/_1129_ ), .ZN(\RegFile/_1130_ ) );
NAND3_X1 \RegFile/_5153_ ( .A1(\RegFile/_0954_ ), .A2(\RegFile/_3738_ ), .A3(\RegFile/_0891_ ), .ZN(\RegFile/_1131_ ) );
AOI22_X1 \RegFile/_5154_ ( .A1(\RegFile/_3770_ ), .A2(\RegFile/_0827_ ), .B1(\RegFile/_0759_ ), .B2(\RegFile/_3642_ ), .ZN(\RegFile/_1132_ ) );
AND4_X1 \RegFile/_5155_ ( .A1(\RegFile/_0814_ ), .A2(\RegFile/_1130_ ), .A3(\RegFile/_1131_ ), .A4(\RegFile/_1132_ ), .ZN(\RegFile/_1133_ ) );
NAND3_X1 \RegFile/_5156_ ( .A1(\RegFile/_0833_ ), .A2(\RegFile/_3354_ ), .A3(\RegFile/_0834_ ), .ZN(\RegFile/_1134_ ) );
INV_X1 \RegFile/_5157_ ( .A(\RegFile/_3578_ ), .ZN(\RegFile/_1135_ ) );
INV_X1 \RegFile/_5158_ ( .A(\RegFile/_3610_ ), .ZN(\RegFile/_1136_ ) );
OAI221_X1 \RegFile/_5159_ ( .A(\RegFile/_1134_ ), .B1(\RegFile/_0838_ ), .B2(\RegFile/_1135_ ), .C1(\RegFile/_0909_ ), .C2(\RegFile/_1136_ ), .ZN(\RegFile/_1137_ ) );
AND3_X1 \RegFile/_5160_ ( .A1(\RegFile/_0841_ ), .A2(\RegFile/_3418_ ), .A3(\RegFile/_0842_ ), .ZN(\RegFile/_1138_ ) );
AND3_X1 \RegFile/_5161_ ( .A1(\RegFile/_0824_ ), .A2(\RegFile/_0784_ ), .A3(\RegFile/_3322_ ), .ZN(\RegFile/_1139_ ) );
NAND3_X1 \RegFile/_5162_ ( .A1(\RegFile/_0765_ ), .A2(\RegFile/_0769_ ), .A3(\RegFile/_3386_ ), .ZN(\RegFile/_1140_ ) );
INV_X1 \RegFile/_5163_ ( .A(\RegFile/_3706_ ), .ZN(\RegFile/_1141_ ) );
OAI21_X1 \RegFile/_5164_ ( .A(\RegFile/_1140_ ), .B1(\RegFile/_0847_ ), .B2(\RegFile/_1141_ ), .ZN(\RegFile/_1142_ ) );
NOR4_X1 \RegFile/_5165_ ( .A1(\RegFile/_1137_ ), .A2(\RegFile/_1138_ ), .A3(\RegFile/_1139_ ), .A4(\RegFile/_1142_ ), .ZN(\RegFile/_1143_ ) );
AOI22_X1 \RegFile/_5166_ ( .A1(\RegFile/_1133_ ), .A2(\RegFile/_1143_ ), .B1(\RegFile/_0080_ ), .B2(\RegFile/_1033_ ), .ZN(\RegFile/_0656_ ) );
NAND3_X1 \RegFile/_5167_ ( .A1(\RegFile/_0943_ ), .A2(\RegFile/_0787_ ), .A3(\RegFile/_3579_ ), .ZN(\RegFile/_1144_ ) );
NAND3_X1 \RegFile/_5168_ ( .A1(\RegFile/_0751_ ), .A2(\RegFile/_0876_ ), .A3(\RegFile/_3323_ ), .ZN(\RegFile/_1145_ ) );
NAND3_X1 \RegFile/_5169_ ( .A1(\RegFile/_0751_ ), .A2(\RegFile/_3355_ ), .A3(\RegFile/_0883_ ), .ZN(\RegFile/_1146_ ) );
NAND2_X1 \RegFile/_5170_ ( .A1(\RegFile/_1145_ ), .A2(\RegFile/_1146_ ), .ZN(\RegFile/_1147_ ) );
AOI221_X4 \RegFile/_5171_ ( .A(\RegFile/_1147_ ), .B1(\RegFile/_3387_ ), .B2(\RegFile/_0872_ ), .C1(\RegFile/_3515_ ), .C2(\RegFile/_0821_ ), .ZN(\RegFile/_1148_ ) );
INV_X1 \RegFile/_5172_ ( .A(\RegFile/_0083_ ), .ZN(\RegFile/_1149_ ) );
AOI22_X1 \RegFile/_5173_ ( .A1(\RegFile/_1149_ ), .A2(\RegFile/_0789_ ), .B1(\RegFile/_0870_ ), .B2(\RegFile/_3611_ ), .ZN(\RegFile/_1150_ ) );
NAND3_X1 \RegFile/_5174_ ( .A1(\RegFile/_0785_ ), .A2(\RegFile/_3547_ ), .A3(\RegFile/_0787_ ), .ZN(\RegFile/_1151_ ) );
AND4_X1 \RegFile/_5175_ ( .A1(\RegFile/_1144_ ), .A2(\RegFile/_1148_ ), .A3(\RegFile/_1150_ ), .A4(\RegFile/_1151_ ), .ZN(\RegFile/_1152_ ) );
NAND3_X1 \RegFile/_5176_ ( .A1(\RegFile/_0841_ ), .A2(\RegFile/_3419_ ), .A3(\RegFile/_0842_ ), .ZN(\RegFile/_1153_ ) );
NAND3_X1 \RegFile/_5177_ ( .A1(\RegFile/_0841_ ), .A2(\RegFile/_0808_ ), .A3(\RegFile/_3643_ ), .ZN(\RegFile/_1154_ ) );
INV_X1 \RegFile/_5178_ ( .A(\RegFile/_3675_ ), .ZN(\RegFile/_1155_ ) );
OAI211_X2 \RegFile/_5179_ ( .A(\RegFile/_1153_ ), .B(\RegFile/_1154_ ), .C1(\RegFile/_0855_ ), .C2(\RegFile/_1155_ ), .ZN(\RegFile/_1156_ ) );
NAND3_X1 \RegFile/_5180_ ( .A1(\RegFile/_0793_ ), .A2(\RegFile/_3739_ ), .A3(\RegFile/_0794_ ), .ZN(\RegFile/_1157_ ) );
INV_X1 \RegFile/_5181_ ( .A(\RegFile/_3707_ ), .ZN(\RegFile/_1158_ ) );
OAI21_X1 \RegFile/_5182_ ( .A(\RegFile/_1157_ ), .B1(\RegFile/_0848_ ), .B2(\RegFile/_1158_ ), .ZN(\RegFile/_1159_ ) );
AND3_X1 \RegFile/_5183_ ( .A1(\RegFile/_0824_ ), .A2(\RegFile/_0796_ ), .A3(\RegFile/_3771_ ), .ZN(\RegFile/_1160_ ) );
NOR4_X1 \RegFile/_5184_ ( .A1(\RegFile/_1156_ ), .A2(\RegFile/_1159_ ), .A3(\RegFile/_0807_ ), .A4(\RegFile/_1160_ ), .ZN(\RegFile/_1161_ ) );
AOI22_X1 \RegFile/_5185_ ( .A1(\RegFile/_1152_ ), .A2(\RegFile/_1161_ ), .B1(\RegFile/_0082_ ), .B2(\RegFile/_1033_ ), .ZN(\RegFile/_0657_ ) );
INV_X1 \RegFile/_5186_ ( .A(\RegFile/_0085_ ), .ZN(\RegFile/_1162_ ) );
AOI22_X1 \RegFile/_5187_ ( .A1(\RegFile/_3644_ ), .A2(\RegFile/_0759_ ), .B1(\RegFile/_0789_ ), .B2(\RegFile/_1162_ ), .ZN(\RegFile/_1163_ ) );
INV_X1 \RegFile/_5188_ ( .A(\RegFile/_3420_ ), .ZN(\RegFile/_1164_ ) );
INV_X1 \RegFile/_5189_ ( .A(\RegFile/_3676_ ), .ZN(\RegFile/_1165_ ) );
OAI221_X1 \RegFile/_5190_ ( .A(\RegFile/_1163_ ), .B1(\RegFile/_1096_ ), .B2(\RegFile/_1164_ ), .C1(\RegFile/_1165_ ), .C2(\RegFile/_0855_ ), .ZN(\RegFile/_1166_ ) );
AND3_X1 \RegFile/_5191_ ( .A1(\RegFile/_0961_ ), .A2(\RegFile/_3356_ ), .A3(\RegFile/_0834_ ), .ZN(\RegFile/_1167_ ) );
AND3_X1 \RegFile/_5192_ ( .A1(\RegFile/_0793_ ), .A2(\RegFile/_0898_ ), .A3(\RegFile/_3324_ ), .ZN(\RegFile/_1168_ ) );
NAND3_X1 \RegFile/_5193_ ( .A1(\RegFile/_0861_ ), .A2(\RegFile/_3516_ ), .A3(\RegFile/_0912_ ), .ZN(\RegFile/_1169_ ) );
NAND3_X1 \RegFile/_5194_ ( .A1(\RegFile/_0842_ ), .A2(\RegFile/_0794_ ), .A3(\RegFile/_3388_ ), .ZN(\RegFile/_1170_ ) );
NAND2_X1 \RegFile/_5195_ ( .A1(\RegFile/_1169_ ), .A2(\RegFile/_1170_ ), .ZN(\RegFile/_1171_ ) );
NOR4_X1 \RegFile/_5196_ ( .A1(\RegFile/_1166_ ), .A2(\RegFile/_1167_ ), .A3(\RegFile/_1168_ ), .A4(\RegFile/_1171_ ), .ZN(\RegFile/_1172_ ) );
NAND3_X1 \RegFile/_5197_ ( .A1(\RegFile/_0898_ ), .A2(\RegFile/_3548_ ), .A3(\RegFile/_0787_ ), .ZN(\RegFile/_1173_ ) );
INV_X1 \RegFile/_5198_ ( .A(\RegFile/_3580_ ), .ZN(\RegFile/_1174_ ) );
INV_X1 \RegFile/_5199_ ( .A(\RegFile/_3612_ ), .ZN(\RegFile/_1175_ ) );
OAI221_X1 \RegFile/_5200_ ( .A(\RegFile/_1173_ ), .B1(\RegFile/_0838_ ), .B2(\RegFile/_1174_ ), .C1(\RegFile/_0909_ ), .C2(\RegFile/_1175_ ), .ZN(\RegFile/_1176_ ) );
NAND3_X1 \RegFile/_5201_ ( .A1(\RegFile/_0824_ ), .A2(\RegFile/_3740_ ), .A3(\RegFile/_0802_ ), .ZN(\RegFile/_1177_ ) );
INV_X1 \RegFile/_5202_ ( .A(\RegFile/_3708_ ), .ZN(\RegFile/_1178_ ) );
OAI21_X1 \RegFile/_5203_ ( .A(\RegFile/_1177_ ), .B1(\RegFile/_0848_ ), .B2(\RegFile/_1178_ ), .ZN(\RegFile/_1179_ ) );
AND3_X1 \RegFile/_5204_ ( .A1(\RegFile/_0824_ ), .A2(\RegFile/_0796_ ), .A3(\RegFile/_3772_ ), .ZN(\RegFile/_1180_ ) );
NOR4_X1 \RegFile/_5205_ ( .A1(\RegFile/_1176_ ), .A2(\RegFile/_0807_ ), .A3(\RegFile/_1179_ ), .A4(\RegFile/_1180_ ), .ZN(\RegFile/_1181_ ) );
AOI22_X1 \RegFile/_5206_ ( .A1(\RegFile/_1172_ ), .A2(\RegFile/_1181_ ), .B1(\RegFile/_0084_ ), .B2(\RegFile/_1033_ ), .ZN(\RegFile/_0658_ ) );
NAND3_X1 \RegFile/_5207_ ( .A1(\RegFile/_0762_ ), .A2(\RegFile/_0897_ ), .A3(\RegFile/_3646_ ), .ZN(\RegFile/_1182_ ) );
INV_X1 \RegFile/_5208_ ( .A(\RegFile/_3678_ ), .ZN(\RegFile/_1183_ ) );
INV_X1 \RegFile/_5209_ ( .A(\RegFile/_3422_ ), .ZN(\RegFile/_1184_ ) );
OAI221_X1 \RegFile/_5210_ ( .A(\RegFile/_1182_ ), .B1(\RegFile/_0855_ ), .B2(\RegFile/_1183_ ), .C1(\RegFile/_1184_ ), .C2(\RegFile/_1096_ ), .ZN(\RegFile/_1185_ ) );
NAND4_X1 \RegFile/_5211_ ( .A1(\RegFile/_0802_ ), .A2(\RegFile/_0643_ ), .A3(\RegFile/_0749_ ), .A4(\RegFile/_3742_ ), .ZN(\RegFile/_1186_ ) );
INV_X1 \RegFile/_5212_ ( .A(\RegFile/_3710_ ), .ZN(\RegFile/_1187_ ) );
OAI21_X1 \RegFile/_5213_ ( .A(\RegFile/_1186_ ), .B1(\RegFile/_0848_ ), .B2(\RegFile/_1187_ ), .ZN(\RegFile/_1188_ ) );
AND3_X1 \RegFile/_5214_ ( .A1(\RegFile/_0844_ ), .A2(\RegFile/_0796_ ), .A3(\RegFile/_3774_ ), .ZN(\RegFile/_1189_ ) );
NOR4_X1 \RegFile/_5215_ ( .A1(\RegFile/_1185_ ), .A2(\RegFile/_0811_ ), .A3(\RegFile/_1188_ ), .A4(\RegFile/_1189_ ), .ZN(\RegFile/_1190_ ) );
AND3_X1 \RegFile/_5216_ ( .A1(\RegFile/_0864_ ), .A2(\RegFile/_3358_ ), .A3(\RegFile/_0775_ ), .ZN(\RegFile/_1191_ ) );
AOI21_X1 \RegFile/_5217_ ( .A(\RegFile/_1191_ ), .B1(\RegFile/_3326_ ), .B2(\RegFile/_0756_ ), .ZN(\RegFile/_1192_ ) );
INV_X1 \RegFile/_5218_ ( .A(\RegFile/_0087_ ), .ZN(\RegFile/_1193_ ) );
AOI22_X1 \RegFile/_5219_ ( .A1(\RegFile/_1193_ ), .A2(\RegFile/_0789_ ), .B1(\RegFile/_0870_ ), .B2(\RegFile/_3614_ ), .ZN(\RegFile/_1194_ ) );
AOI22_X1 \RegFile/_5220_ ( .A1(\RegFile/_0822_ ), .A2(\RegFile/_3518_ ), .B1(\RegFile/_0872_ ), .B2(\RegFile/_3390_ ), .ZN(\RegFile/_1195_ ) );
AOI22_X1 \RegFile/_5221_ ( .A1(\RegFile/_0820_ ), .A2(\RegFile/_3550_ ), .B1(\RegFile/_0780_ ), .B2(\RegFile/_3582_ ), .ZN(\RegFile/_1196_ ) );
AND4_X1 \RegFile/_5222_ ( .A1(\RegFile/_1192_ ), .A2(\RegFile/_1194_ ), .A3(\RegFile/_1195_ ), .A4(\RegFile/_1196_ ), .ZN(\RegFile/_1197_ ) );
BUF_X4 \RegFile/_5223_ ( .A(\RegFile/_0807_ ), .Z(\RegFile/_1198_ ) );
AOI22_X1 \RegFile/_5224_ ( .A1(\RegFile/_1190_ ), .A2(\RegFile/_1197_ ), .B1(\RegFile/_0086_ ), .B2(\RegFile/_1198_ ), .ZN(\RegFile/_0660_ ) );
AND3_X1 \RegFile/_5225_ ( .A1(\RegFile/_0751_ ), .A2(\RegFile/_3359_ ), .A3(\RegFile/_0774_ ), .ZN(\RegFile/_1199_ ) );
AOI221_X4 \RegFile/_5226_ ( .A(\RegFile/_1199_ ), .B1(\RegFile/_3583_ ), .B2(\RegFile/_0779_ ), .C1(\RegFile/_3615_ ), .C2(\RegFile/_0870_ ), .ZN(\RegFile/_1200_ ) );
AND3_X1 \RegFile/_5227_ ( .A1(\RegFile/_0864_ ), .A2(\RegFile/_0949_ ), .A3(\RegFile/_3327_ ), .ZN(\RegFile/_1201_ ) );
AOI21_X1 \RegFile/_5228_ ( .A(\RegFile/_1201_ ), .B1(\RegFile/_3423_ ), .B2(\RegFile/_0889_ ), .ZN(\RegFile/_1202_ ) );
NAND3_X1 \RegFile/_5229_ ( .A1(\RegFile/_0766_ ), .A2(\RegFile/_0770_ ), .A3(\RegFile/_3391_ ), .ZN(\RegFile/_1203_ ) );
NAND3_X1 \RegFile/_5230_ ( .A1(\RegFile/_0893_ ), .A2(\RegFile/_3711_ ), .A3(\RegFile/_0943_ ), .ZN(\RegFile/_1204_ ) );
AND4_X1 \RegFile/_5231_ ( .A1(\RegFile/_1200_ ), .A2(\RegFile/_1202_ ), .A3(\RegFile/_1203_ ), .A4(\RegFile/_1204_ ), .ZN(\RegFile/_1205_ ) );
AOI22_X1 \RegFile/_5232_ ( .A1(\RegFile/_3775_ ), .A2(\RegFile/_0828_ ), .B1(\RegFile/_0829_ ), .B2(\RegFile/_3647_ ), .ZN(\RegFile/_1206_ ) );
NAND3_X1 \RegFile/_5233_ ( .A1(\RegFile/_0761_ ), .A2(\RegFile/_3519_ ), .A3(\RegFile/_0786_ ), .ZN(\RegFile/_1207_ ) );
NAND3_X1 \RegFile/_5234_ ( .A1(\RegFile/_0801_ ), .A2(\RegFile/_0886_ ), .A3(\RegFile/_3679_ ), .ZN(\RegFile/_1208_ ) );
NAND3_X1 \RegFile/_5235_ ( .A1(\RegFile/_0949_ ), .A2(\RegFile/_3551_ ), .A3(\RegFile/_0786_ ), .ZN(\RegFile/_1209_ ) );
INV_X1 \RegFile/_5236_ ( .A(\RegFile/_0089_ ), .ZN(\RegFile/_1210_ ) );
NAND3_X1 \RegFile/_5237_ ( .A1(\RegFile/_0783_ ), .A2(\RegFile/_1210_ ), .A3(\RegFile/_0764_ ), .ZN(\RegFile/_1211_ ) );
AND4_X1 \RegFile/_5238_ ( .A1(\RegFile/_1207_ ), .A2(\RegFile/_1208_ ), .A3(\RegFile/_1209_ ), .A4(\RegFile/_1211_ ), .ZN(\RegFile/_1212_ ) );
NAND3_X1 \RegFile/_5239_ ( .A1(\RegFile/_0954_ ), .A2(\RegFile/_3743_ ), .A3(\RegFile/_0955_ ), .ZN(\RegFile/_1213_ ) );
AND4_X1 \RegFile/_5240_ ( .A1(\RegFile/_0813_ ), .A2(\RegFile/_1206_ ), .A3(\RegFile/_1212_ ), .A4(\RegFile/_1213_ ), .ZN(\RegFile/_1214_ ) );
AOI22_X1 \RegFile/_5241_ ( .A1(\RegFile/_1205_ ), .A2(\RegFile/_1214_ ), .B1(\RegFile/_0088_ ), .B2(\RegFile/_1198_ ), .ZN(\RegFile/_0661_ ) );
AND3_X1 \RegFile/_5242_ ( .A1(\RegFile/_0751_ ), .A2(\RegFile/_3360_ ), .A3(\RegFile/_0883_ ), .ZN(\RegFile/_1215_ ) );
AOI221_X4 \RegFile/_5243_ ( .A(\RegFile/_1215_ ), .B1(\RegFile/_3584_ ), .B2(\RegFile/_0779_ ), .C1(\RegFile/_3616_ ), .C2(\RegFile/_0870_ ), .ZN(\RegFile/_1216_ ) );
AND3_X1 \RegFile/_5244_ ( .A1(\RegFile/_0832_ ), .A2(\RegFile/_0949_ ), .A3(\RegFile/_3328_ ), .ZN(\RegFile/_1217_ ) );
AOI21_X1 \RegFile/_5245_ ( .A(\RegFile/_1217_ ), .B1(\RegFile/_3424_ ), .B2(\RegFile/_0889_ ), .ZN(\RegFile/_1218_ ) );
NAND3_X1 \RegFile/_5246_ ( .A1(\RegFile/_0766_ ), .A2(\RegFile/_0770_ ), .A3(\RegFile/_3392_ ), .ZN(\RegFile/_1219_ ) );
NAND3_X1 \RegFile/_5247_ ( .A1(\RegFile/_0893_ ), .A2(\RegFile/_3712_ ), .A3(\RegFile/_0943_ ), .ZN(\RegFile/_1220_ ) );
AND4_X1 \RegFile/_5248_ ( .A1(\RegFile/_1216_ ), .A2(\RegFile/_1218_ ), .A3(\RegFile/_1219_ ), .A4(\RegFile/_1220_ ), .ZN(\RegFile/_1221_ ) );
AOI22_X1 \RegFile/_5249_ ( .A1(\RegFile/_3776_ ), .A2(\RegFile/_0828_ ), .B1(\RegFile/_0829_ ), .B2(\RegFile/_3648_ ), .ZN(\RegFile/_1222_ ) );
NAND3_X1 \RegFile/_5250_ ( .A1(\RegFile/_0761_ ), .A2(\RegFile/_3520_ ), .A3(\RegFile/_0786_ ), .ZN(\RegFile/_1223_ ) );
NAND3_X1 \RegFile/_5251_ ( .A1(\RegFile/_0800_ ), .A2(\RegFile/_0886_ ), .A3(\RegFile/_3680_ ), .ZN(\RegFile/_1224_ ) );
NAND3_X1 \RegFile/_5252_ ( .A1(\RegFile/_0949_ ), .A2(\RegFile/_3552_ ), .A3(\RegFile/_0786_ ), .ZN(\RegFile/_1225_ ) );
INV_X1 \RegFile/_5253_ ( .A(\RegFile/_0091_ ), .ZN(\RegFile/_1226_ ) );
NAND3_X1 \RegFile/_5254_ ( .A1(\RegFile/_0783_ ), .A2(\RegFile/_1226_ ), .A3(\RegFile/_0764_ ), .ZN(\RegFile/_1227_ ) );
AND4_X1 \RegFile/_5255_ ( .A1(\RegFile/_1223_ ), .A2(\RegFile/_1224_ ), .A3(\RegFile/_1225_ ), .A4(\RegFile/_1227_ ), .ZN(\RegFile/_1228_ ) );
NAND3_X1 \RegFile/_5256_ ( .A1(\RegFile/_0961_ ), .A2(\RegFile/_3744_ ), .A3(\RegFile/_0955_ ), .ZN(\RegFile/_1229_ ) );
AND4_X1 \RegFile/_5257_ ( .A1(\RegFile/_0813_ ), .A2(\RegFile/_1222_ ), .A3(\RegFile/_1228_ ), .A4(\RegFile/_1229_ ), .ZN(\RegFile/_1230_ ) );
AOI22_X1 \RegFile/_5258_ ( .A1(\RegFile/_1221_ ), .A2(\RegFile/_1230_ ), .B1(\RegFile/_0090_ ), .B2(\RegFile/_1198_ ), .ZN(\RegFile/_0662_ ) );
AND3_X1 \RegFile/_5259_ ( .A1(\RegFile/_0751_ ), .A2(\RegFile/_3361_ ), .A3(\RegFile/_0883_ ), .ZN(\RegFile/_1231_ ) );
AOI221_X4 \RegFile/_5260_ ( .A(\RegFile/_1231_ ), .B1(\RegFile/_3617_ ), .B2(\RegFile/_0869_ ), .C1(\RegFile/_3585_ ), .C2(\RegFile/_0780_ ), .ZN(\RegFile/_1232_ ) );
AND3_X1 \RegFile/_5261_ ( .A1(\RegFile/_0832_ ), .A2(\RegFile/_0949_ ), .A3(\RegFile/_3329_ ), .ZN(\RegFile/_1233_ ) );
AOI21_X1 \RegFile/_5262_ ( .A(\RegFile/_1233_ ), .B1(\RegFile/_3425_ ), .B2(\RegFile/_0889_ ), .ZN(\RegFile/_1234_ ) );
NAND3_X1 \RegFile/_5263_ ( .A1(\RegFile/_0766_ ), .A2(\RegFile/_0770_ ), .A3(\RegFile/_3393_ ), .ZN(\RegFile/_1235_ ) );
NAND3_X1 \RegFile/_5264_ ( .A1(\RegFile/_0893_ ), .A2(\RegFile/_3713_ ), .A3(\RegFile/_0943_ ), .ZN(\RegFile/_1236_ ) );
AND4_X1 \RegFile/_5265_ ( .A1(\RegFile/_1232_ ), .A2(\RegFile/_1234_ ), .A3(\RegFile/_1235_ ), .A4(\RegFile/_1236_ ), .ZN(\RegFile/_1237_ ) );
AOI22_X1 \RegFile/_5266_ ( .A1(\RegFile/_3777_ ), .A2(\RegFile/_0828_ ), .B1(\RegFile/_0829_ ), .B2(\RegFile/_3649_ ), .ZN(\RegFile/_1238_ ) );
NAND3_X1 \RegFile/_5267_ ( .A1(\RegFile/_0761_ ), .A2(\RegFile/_3521_ ), .A3(\RegFile/_0786_ ), .ZN(\RegFile/_1239_ ) );
NAND3_X1 \RegFile/_5268_ ( .A1(\RegFile/_0800_ ), .A2(\RegFile/_0886_ ), .A3(\RegFile/_3681_ ), .ZN(\RegFile/_1240_ ) );
NAND3_X1 \RegFile/_5269_ ( .A1(\RegFile/_0949_ ), .A2(\RegFile/_3553_ ), .A3(\RegFile/_0777_ ), .ZN(\RegFile/_1241_ ) );
INV_X1 \RegFile/_5270_ ( .A(\RegFile/_0093_ ), .ZN(\RegFile/_1242_ ) );
NAND3_X1 \RegFile/_5271_ ( .A1(\RegFile/_0783_ ), .A2(\RegFile/_1242_ ), .A3(\RegFile/_0764_ ), .ZN(\RegFile/_1243_ ) );
AND4_X1 \RegFile/_5272_ ( .A1(\RegFile/_1239_ ), .A2(\RegFile/_1240_ ), .A3(\RegFile/_1241_ ), .A4(\RegFile/_1243_ ), .ZN(\RegFile/_1244_ ) );
NAND3_X1 \RegFile/_5273_ ( .A1(\RegFile/_0961_ ), .A2(\RegFile/_3745_ ), .A3(\RegFile/_0955_ ), .ZN(\RegFile/_1245_ ) );
AND4_X1 \RegFile/_5274_ ( .A1(\RegFile/_0813_ ), .A2(\RegFile/_1238_ ), .A3(\RegFile/_1244_ ), .A4(\RegFile/_1245_ ), .ZN(\RegFile/_1246_ ) );
AOI22_X1 \RegFile/_5275_ ( .A1(\RegFile/_1237_ ), .A2(\RegFile/_1246_ ), .B1(\RegFile/_0092_ ), .B2(\RegFile/_1198_ ), .ZN(\RegFile/_0663_ ) );
NAND3_X1 \RegFile/_5276_ ( .A1(\RegFile/_0762_ ), .A2(\RegFile/_0808_ ), .A3(\RegFile/_3650_ ), .ZN(\RegFile/_1247_ ) );
INV_X1 \RegFile/_5277_ ( .A(\RegFile/_3682_ ), .ZN(\RegFile/_1248_ ) );
INV_X1 \RegFile/_5278_ ( .A(\RegFile/_3426_ ), .ZN(\RegFile/_1249_ ) );
OAI221_X1 \RegFile/_5279_ ( .A(\RegFile/_1247_ ), .B1(\RegFile/_0855_ ), .B2(\RegFile/_1248_ ), .C1(\RegFile/_1249_ ), .C2(\RegFile/_1096_ ), .ZN(\RegFile/_1250_ ) );
NAND3_X1 \RegFile/_5280_ ( .A1(\RegFile/_0833_ ), .A2(\RegFile/_3746_ ), .A3(\RegFile/_0836_ ), .ZN(\RegFile/_1251_ ) );
NAND3_X1 \RegFile/_5281_ ( .A1(\RegFile/_0808_ ), .A2(\RegFile/_3714_ ), .A3(\RegFile/_0918_ ), .ZN(\RegFile/_1252_ ) );
NAND2_X1 \RegFile/_5282_ ( .A1(\RegFile/_1251_ ), .A2(\RegFile/_1252_ ), .ZN(\RegFile/_1253_ ) );
AND3_X1 \RegFile/_5283_ ( .A1(\RegFile/_0844_ ), .A2(\RegFile/_0796_ ), .A3(\RegFile/_3778_ ), .ZN(\RegFile/_1254_ ) );
NOR4_X1 \RegFile/_5284_ ( .A1(\RegFile/_1250_ ), .A2(\RegFile/_0811_ ), .A3(\RegFile/_1253_ ), .A4(\RegFile/_1254_ ), .ZN(\RegFile/_1255_ ) );
AND3_X1 \RegFile/_5285_ ( .A1(\RegFile/_0864_ ), .A2(\RegFile/_3362_ ), .A3(\RegFile/_0775_ ), .ZN(\RegFile/_1256_ ) );
AOI21_X1 \RegFile/_5286_ ( .A(\RegFile/_1256_ ), .B1(\RegFile/_3330_ ), .B2(\RegFile/_0756_ ), .ZN(\RegFile/_1257_ ) );
INV_X1 \RegFile/_5287_ ( .A(\RegFile/_0095_ ), .ZN(\RegFile/_1258_ ) );
AOI22_X1 \RegFile/_5288_ ( .A1(\RegFile/_1258_ ), .A2(\RegFile/_0789_ ), .B1(\RegFile/_0870_ ), .B2(\RegFile/_3618_ ), .ZN(\RegFile/_1259_ ) );
AOI22_X1 \RegFile/_5289_ ( .A1(\RegFile/_0822_ ), .A2(\RegFile/_3522_ ), .B1(\RegFile/_0872_ ), .B2(\RegFile/_3394_ ), .ZN(\RegFile/_1260_ ) );
AOI22_X1 \RegFile/_5290_ ( .A1(\RegFile/_0820_ ), .A2(\RegFile/_3554_ ), .B1(\RegFile/_0780_ ), .B2(\RegFile/_3586_ ), .ZN(\RegFile/_1261_ ) );
AND4_X1 \RegFile/_5291_ ( .A1(\RegFile/_1257_ ), .A2(\RegFile/_1259_ ), .A3(\RegFile/_1260_ ), .A4(\RegFile/_1261_ ), .ZN(\RegFile/_1262_ ) );
AOI22_X1 \RegFile/_5292_ ( .A1(\RegFile/_1255_ ), .A2(\RegFile/_1262_ ), .B1(\RegFile/_0094_ ), .B2(\RegFile/_1198_ ), .ZN(\RegFile/_0664_ ) );
NAND3_X1 \RegFile/_5293_ ( .A1(\RegFile/_0825_ ), .A2(\RegFile/_3363_ ), .A3(\RegFile/_0943_ ), .ZN(\RegFile/_1263_ ) );
INV_X1 \RegFile/_5294_ ( .A(\RegFile/_3651_ ), .ZN(\RegFile/_1264_ ) );
OAI22_X1 \RegFile/_5295_ ( .A1(\RegFile/_0901_ ), .A2(\RegFile/_1264_ ), .B1(\RegFile/_0790_ ), .B2(\RegFile/_0097_ ), .ZN(\RegFile/_1265_ ) );
AOI221_X4 \RegFile/_5296_ ( .A(\RegFile/_1265_ ), .B1(\RegFile/_3427_ ), .B2(\RegFile/_0888_ ), .C1(\RegFile/_3683_ ), .C2(\RegFile/_0815_ ), .ZN(\RegFile/_1266_ ) );
NAND3_X1 \RegFile/_5297_ ( .A1(\RegFile/_0954_ ), .A2(\RegFile/_0785_ ), .A3(\RegFile/_3331_ ), .ZN(\RegFile/_1267_ ) );
AOI22_X1 \RegFile/_5298_ ( .A1(\RegFile/_0822_ ), .A2(\RegFile/_3523_ ), .B1(\RegFile/_0872_ ), .B2(\RegFile/_3395_ ), .ZN(\RegFile/_1268_ ) );
AND4_X1 \RegFile/_5299_ ( .A1(\RegFile/_1263_ ), .A2(\RegFile/_1266_ ), .A3(\RegFile/_1267_ ), .A4(\RegFile/_1268_ ), .ZN(\RegFile/_1269_ ) );
NAND3_X1 \RegFile/_5300_ ( .A1(\RegFile/_0808_ ), .A2(\RegFile/_3619_ ), .A3(\RegFile/_0836_ ), .ZN(\RegFile/_1270_ ) );
INV_X1 \RegFile/_5301_ ( .A(\RegFile/_3587_ ), .ZN(\RegFile/_1271_ ) );
INV_X1 \RegFile/_5302_ ( .A(\RegFile/_3555_ ), .ZN(\RegFile/_1272_ ) );
OAI221_X1 \RegFile/_5303_ ( .A(\RegFile/_1270_ ), .B1(\RegFile/_0838_ ), .B2(\RegFile/_1271_ ), .C1(\RegFile/_0914_ ), .C2(\RegFile/_1272_ ), .ZN(\RegFile/_1273_ ) );
NAND3_X1 \RegFile/_5304_ ( .A1(\RegFile/_0824_ ), .A2(\RegFile/_3747_ ), .A3(\RegFile/_0802_ ), .ZN(\RegFile/_1274_ ) );
INV_X1 \RegFile/_5305_ ( .A(\RegFile/_3715_ ), .ZN(\RegFile/_1275_ ) );
OAI21_X1 \RegFile/_5306_ ( .A(\RegFile/_1274_ ), .B1(\RegFile/_0848_ ), .B2(\RegFile/_1275_ ), .ZN(\RegFile/_1276_ ) );
AND3_X1 \RegFile/_5307_ ( .A1(\RegFile/_0824_ ), .A2(\RegFile/_0796_ ), .A3(\RegFile/_3779_ ), .ZN(\RegFile/_1277_ ) );
NOR4_X1 \RegFile/_5308_ ( .A1(\RegFile/_1273_ ), .A2(\RegFile/_0807_ ), .A3(\RegFile/_1276_ ), .A4(\RegFile/_1277_ ), .ZN(\RegFile/_1278_ ) );
AOI22_X1 \RegFile/_5309_ ( .A1(\RegFile/_1269_ ), .A2(\RegFile/_1278_ ), .B1(\RegFile/_0096_ ), .B2(\RegFile/_1198_ ), .ZN(\RegFile/_0665_ ) );
NAND3_X1 \RegFile/_5310_ ( .A1(\RegFile/_0762_ ), .A2(\RegFile/_3428_ ), .A3(\RegFile/_0852_ ), .ZN(\RegFile/_1279_ ) );
INV_X1 \RegFile/_5311_ ( .A(\RegFile/_3684_ ), .ZN(\RegFile/_1280_ ) );
INV_X1 \RegFile/_5312_ ( .A(\RegFile/_3652_ ), .ZN(\RegFile/_1281_ ) );
OAI221_X1 \RegFile/_5313_ ( .A(\RegFile/_1279_ ), .B1(\RegFile/_0855_ ), .B2(\RegFile/_1280_ ), .C1(\RegFile/_1281_ ), .C2(\RegFile/_0901_ ), .ZN(\RegFile/_1282_ ) );
NAND3_X1 \RegFile/_5314_ ( .A1(\RegFile/_0833_ ), .A2(\RegFile/_3748_ ), .A3(\RegFile/_0836_ ), .ZN(\RegFile/_1283_ ) );
NAND3_X1 \RegFile/_5315_ ( .A1(\RegFile/_0808_ ), .A2(\RegFile/_3716_ ), .A3(\RegFile/_0918_ ), .ZN(\RegFile/_1284_ ) );
NAND2_X1 \RegFile/_5316_ ( .A1(\RegFile/_1283_ ), .A2(\RegFile/_1284_ ), .ZN(\RegFile/_1285_ ) );
AND3_X1 \RegFile/_5317_ ( .A1(\RegFile/_0844_ ), .A2(\RegFile/_0796_ ), .A3(\RegFile/_3780_ ), .ZN(\RegFile/_1286_ ) );
NOR4_X1 \RegFile/_5318_ ( .A1(\RegFile/_1282_ ), .A2(\RegFile/_0811_ ), .A3(\RegFile/_1285_ ), .A4(\RegFile/_1286_ ), .ZN(\RegFile/_1287_ ) );
NAND3_X1 \RegFile/_5319_ ( .A1(\RegFile/_0897_ ), .A2(\RegFile/_3620_ ), .A3(\RegFile/_0836_ ), .ZN(\RegFile/_1288_ ) );
OAI21_X1 \RegFile/_5320_ ( .A(\RegFile/_1288_ ), .B1(\RegFile/_0791_ ), .B2(\RegFile/_0099_ ), .ZN(\RegFile/_1289_ ) );
NAND3_X1 \RegFile/_5321_ ( .A1(\RegFile/_0961_ ), .A2(\RegFile/_0785_ ), .A3(\RegFile/_3332_ ), .ZN(\RegFile/_1290_ ) );
NAND3_X1 \RegFile/_5322_ ( .A1(\RegFile/_0833_ ), .A2(\RegFile/_3364_ ), .A3(\RegFile/_0834_ ), .ZN(\RegFile/_1291_ ) );
NAND2_X1 \RegFile/_5323_ ( .A1(\RegFile/_1290_ ), .A2(\RegFile/_1291_ ), .ZN(\RegFile/_1292_ ) );
NAND3_X1 \RegFile/_5324_ ( .A1(\RegFile/_0861_ ), .A2(\RegFile/_3524_ ), .A3(\RegFile/_0912_ ), .ZN(\RegFile/_1293_ ) );
NAND3_X1 \RegFile/_5325_ ( .A1(\RegFile/_0842_ ), .A2(\RegFile/_0794_ ), .A3(\RegFile/_3396_ ), .ZN(\RegFile/_1294_ ) );
NAND2_X1 \RegFile/_5326_ ( .A1(\RegFile/_1293_ ), .A2(\RegFile/_1294_ ), .ZN(\RegFile/_1295_ ) );
NAND3_X1 \RegFile/_5327_ ( .A1(\RegFile/_0898_ ), .A2(\RegFile/_3556_ ), .A3(\RegFile/_0797_ ), .ZN(\RegFile/_1296_ ) );
NAND3_X1 \RegFile/_5328_ ( .A1(\RegFile/_0918_ ), .A2(\RegFile/_0797_ ), .A3(\RegFile/_3588_ ), .ZN(\RegFile/_1297_ ) );
NAND2_X1 \RegFile/_5329_ ( .A1(\RegFile/_1296_ ), .A2(\RegFile/_1297_ ), .ZN(\RegFile/_1298_ ) );
NOR4_X1 \RegFile/_5330_ ( .A1(\RegFile/_1289_ ), .A2(\RegFile/_1292_ ), .A3(\RegFile/_1295_ ), .A4(\RegFile/_1298_ ), .ZN(\RegFile/_1299_ ) );
AOI22_X1 \RegFile/_5331_ ( .A1(\RegFile/_1287_ ), .A2(\RegFile/_1299_ ), .B1(\RegFile/_0098_ ), .B2(\RegFile/_1198_ ), .ZN(\RegFile/_0666_ ) );
NAND3_X1 \RegFile/_5332_ ( .A1(\RegFile/_0799_ ), .A2(\RegFile/_0876_ ), .A3(\RegFile/_3685_ ), .ZN(\RegFile/_1300_ ) );
OAI21_X1 \RegFile/_5333_ ( .A(\RegFile/_1300_ ), .B1(\RegFile/_0790_ ), .B2(\RegFile/_0101_ ), .ZN(\RegFile/_1301_ ) );
AOI221_X4 \RegFile/_5334_ ( .A(\RegFile/_1301_ ), .B1(\RegFile/_3557_ ), .B2(\RegFile/_0819_ ), .C1(\RegFile/_3525_ ), .C2(\RegFile/_0821_ ), .ZN(\RegFile/_1302_ ) );
NAND3_X1 \RegFile/_5335_ ( .A1(\RegFile/_0954_ ), .A2(\RegFile/_3749_ ), .A3(\RegFile/_0891_ ), .ZN(\RegFile/_1303_ ) );
AOI22_X1 \RegFile/_5336_ ( .A1(\RegFile/_3781_ ), .A2(\RegFile/_0827_ ), .B1(\RegFile/_0759_ ), .B2(\RegFile/_3653_ ), .ZN(\RegFile/_1304_ ) );
AND4_X1 \RegFile/_5337_ ( .A1(\RegFile/_0814_ ), .A2(\RegFile/_1302_ ), .A3(\RegFile/_1303_ ), .A4(\RegFile/_1304_ ), .ZN(\RegFile/_1305_ ) );
AND3_X1 \RegFile/_5338_ ( .A1(\RegFile/_0750_ ), .A2(\RegFile/_3365_ ), .A3(\RegFile/_0883_ ), .ZN(\RegFile/_1306_ ) );
AOI221_X4 \RegFile/_5339_ ( .A(\RegFile/_1306_ ), .B1(\RegFile/_3621_ ), .B2(\RegFile/_0869_ ), .C1(\RegFile/_3589_ ), .C2(\RegFile/_0779_ ), .ZN(\RegFile/_1307_ ) );
AND3_X1 \RegFile/_5340_ ( .A1(\RegFile/_0772_ ), .A2(\RegFile/_0783_ ), .A3(\RegFile/_3333_ ), .ZN(\RegFile/_1308_ ) );
AOI21_X1 \RegFile/_5341_ ( .A(\RegFile/_1308_ ), .B1(\RegFile/_3429_ ), .B2(\RegFile/_0888_ ), .ZN(\RegFile/_1309_ ) );
NAND3_X1 \RegFile/_5342_ ( .A1(\RegFile/_0852_ ), .A2(\RegFile/_0955_ ), .A3(\RegFile/_3397_ ), .ZN(\RegFile/_1310_ ) );
NAND3_X1 \RegFile/_5343_ ( .A1(\RegFile/_0897_ ), .A2(\RegFile/_3717_ ), .A3(\RegFile/_0894_ ), .ZN(\RegFile/_1311_ ) );
AND4_X1 \RegFile/_5344_ ( .A1(\RegFile/_1307_ ), .A2(\RegFile/_1309_ ), .A3(\RegFile/_1310_ ), .A4(\RegFile/_1311_ ), .ZN(\RegFile/_1312_ ) );
AOI22_X1 \RegFile/_5345_ ( .A1(\RegFile/_1305_ ), .A2(\RegFile/_1312_ ), .B1(\RegFile/_0100_ ), .B2(\RegFile/_1198_ ), .ZN(\RegFile/_0667_ ) );
NAND3_X1 \RegFile/_5346_ ( .A1(\RegFile/_0762_ ), .A2(\RegFile/_3430_ ), .A3(\RegFile/_0852_ ), .ZN(\RegFile/_1313_ ) );
INV_X1 \RegFile/_5347_ ( .A(\RegFile/_3686_ ), .ZN(\RegFile/_1314_ ) );
INV_X1 \RegFile/_5348_ ( .A(\RegFile/_3654_ ), .ZN(\RegFile/_1315_ ) );
OAI221_X1 \RegFile/_5349_ ( .A(\RegFile/_1313_ ), .B1(\RegFile/_0855_ ), .B2(\RegFile/_1314_ ), .C1(\RegFile/_1315_ ), .C2(\RegFile/_0901_ ), .ZN(\RegFile/_1316_ ) );
NAND4_X1 \RegFile/_5350_ ( .A1(\RegFile/_0802_ ), .A2(\RegFile/_0643_ ), .A3(\RegFile/_0749_ ), .A4(\RegFile/_3750_ ), .ZN(\RegFile/_1317_ ) );
INV_X1 \RegFile/_5351_ ( .A(\RegFile/_3718_ ), .ZN(\RegFile/_1318_ ) );
OAI21_X1 \RegFile/_5352_ ( .A(\RegFile/_1317_ ), .B1(\RegFile/_0848_ ), .B2(\RegFile/_1318_ ), .ZN(\RegFile/_1319_ ) );
AND3_X1 \RegFile/_5353_ ( .A1(\RegFile/_0844_ ), .A2(\RegFile/_0796_ ), .A3(\RegFile/_3782_ ), .ZN(\RegFile/_1320_ ) );
NOR4_X1 \RegFile/_5354_ ( .A1(\RegFile/_1316_ ), .A2(\RegFile/_0811_ ), .A3(\RegFile/_1319_ ), .A4(\RegFile/_1320_ ), .ZN(\RegFile/_1321_ ) );
AND3_X1 \RegFile/_5355_ ( .A1(\RegFile/_0824_ ), .A2(\RegFile/_3366_ ), .A3(\RegFile/_0775_ ), .ZN(\RegFile/_1322_ ) );
AND3_X1 \RegFile/_5356_ ( .A1(\RegFile/_0864_ ), .A2(\RegFile/_0784_ ), .A3(\RegFile/_3334_ ), .ZN(\RegFile/_1323_ ) );
OR2_X1 \RegFile/_5357_ ( .A1(\RegFile/_1322_ ), .A2(\RegFile/_1323_ ), .ZN(\RegFile/_1324_ ) );
NAND3_X1 \RegFile/_5358_ ( .A1(\RegFile/_0808_ ), .A2(\RegFile/_3622_ ), .A3(\RegFile/_0794_ ), .ZN(\RegFile/_1325_ ) );
OAI21_X1 \RegFile/_5359_ ( .A(\RegFile/_1325_ ), .B1(\RegFile/_0791_ ), .B2(\RegFile/_0103_ ), .ZN(\RegFile/_1326_ ) );
NAND3_X1 \RegFile/_5360_ ( .A1(\RegFile/_0861_ ), .A2(\RegFile/_3526_ ), .A3(\RegFile/_0912_ ), .ZN(\RegFile/_1327_ ) );
NAND3_X1 \RegFile/_5361_ ( .A1(\RegFile/_0765_ ), .A2(\RegFile/_0794_ ), .A3(\RegFile/_3398_ ), .ZN(\RegFile/_1328_ ) );
NAND2_X1 \RegFile/_5362_ ( .A1(\RegFile/_1327_ ), .A2(\RegFile/_1328_ ), .ZN(\RegFile/_1329_ ) );
NAND3_X1 \RegFile/_5363_ ( .A1(\RegFile/_0898_ ), .A2(\RegFile/_3558_ ), .A3(\RegFile/_0797_ ), .ZN(\RegFile/_1330_ ) );
NAND3_X1 \RegFile/_5364_ ( .A1(\RegFile/_0918_ ), .A2(\RegFile/_0797_ ), .A3(\RegFile/_3590_ ), .ZN(\RegFile/_1331_ ) );
NAND2_X1 \RegFile/_5365_ ( .A1(\RegFile/_1330_ ), .A2(\RegFile/_1331_ ), .ZN(\RegFile/_1332_ ) );
NOR4_X1 \RegFile/_5366_ ( .A1(\RegFile/_1324_ ), .A2(\RegFile/_1326_ ), .A3(\RegFile/_1329_ ), .A4(\RegFile/_1332_ ), .ZN(\RegFile/_1333_ ) );
AOI22_X1 \RegFile/_5367_ ( .A1(\RegFile/_1321_ ), .A2(\RegFile/_1333_ ), .B1(\RegFile/_0102_ ), .B2(\RegFile/_1198_ ), .ZN(\RegFile/_0668_ ) );
AND3_X1 \RegFile/_5368_ ( .A1(\RegFile/_0751_ ), .A2(\RegFile/_3367_ ), .A3(\RegFile/_0883_ ), .ZN(\RegFile/_1334_ ) );
AOI221_X4 \RegFile/_5369_ ( .A(\RegFile/_1334_ ), .B1(\RegFile/_3623_ ), .B2(\RegFile/_0869_ ), .C1(\RegFile/_3591_ ), .C2(\RegFile/_0780_ ), .ZN(\RegFile/_1335_ ) );
AND3_X1 \RegFile/_5370_ ( .A1(\RegFile/_0832_ ), .A2(\RegFile/_0949_ ), .A3(\RegFile/_3335_ ), .ZN(\RegFile/_1336_ ) );
AOI21_X1 \RegFile/_5371_ ( .A(\RegFile/_1336_ ), .B1(\RegFile/_3431_ ), .B2(\RegFile/_0889_ ), .ZN(\RegFile/_1337_ ) );
NAND3_X1 \RegFile/_5372_ ( .A1(\RegFile/_0766_ ), .A2(\RegFile/_0770_ ), .A3(\RegFile/_3399_ ), .ZN(\RegFile/_1338_ ) );
NAND3_X1 \RegFile/_5373_ ( .A1(\RegFile/_0893_ ), .A2(\RegFile/_3719_ ), .A3(\RegFile/_0894_ ), .ZN(\RegFile/_1339_ ) );
AND4_X1 \RegFile/_5374_ ( .A1(\RegFile/_1335_ ), .A2(\RegFile/_1337_ ), .A3(\RegFile/_1338_ ), .A4(\RegFile/_1339_ ), .ZN(\RegFile/_1340_ ) );
AOI22_X1 \RegFile/_5375_ ( .A1(\RegFile/_3783_ ), .A2(\RegFile/_0828_ ), .B1(\RegFile/_0829_ ), .B2(\RegFile/_3655_ ), .ZN(\RegFile/_1341_ ) );
NAND3_X1 \RegFile/_5376_ ( .A1(\RegFile/_0761_ ), .A2(\RegFile/_3527_ ), .A3(\RegFile/_0786_ ), .ZN(\RegFile/_1342_ ) );
NAND3_X1 \RegFile/_5377_ ( .A1(\RegFile/_0800_ ), .A2(\RegFile/_0886_ ), .A3(\RegFile/_3687_ ), .ZN(\RegFile/_1343_ ) );
NAND3_X1 \RegFile/_5378_ ( .A1(\RegFile/_0949_ ), .A2(\RegFile/_3559_ ), .A3(\RegFile/_0777_ ), .ZN(\RegFile/_1344_ ) );
INV_X1 \RegFile/_5379_ ( .A(\RegFile/_0105_ ), .ZN(\RegFile/_1345_ ) );
NAND3_X1 \RegFile/_5380_ ( .A1(\RegFile/_0783_ ), .A2(\RegFile/_1345_ ), .A3(\RegFile/_0764_ ), .ZN(\RegFile/_1346_ ) );
AND4_X1 \RegFile/_5381_ ( .A1(\RegFile/_1342_ ), .A2(\RegFile/_1343_ ), .A3(\RegFile/_1344_ ), .A4(\RegFile/_1346_ ), .ZN(\RegFile/_1347_ ) );
NAND3_X1 \RegFile/_5382_ ( .A1(\RegFile/_0961_ ), .A2(\RegFile/_3751_ ), .A3(\RegFile/_0955_ ), .ZN(\RegFile/_1348_ ) );
AND4_X1 \RegFile/_5383_ ( .A1(\RegFile/_0813_ ), .A2(\RegFile/_1341_ ), .A3(\RegFile/_1347_ ), .A4(\RegFile/_1348_ ), .ZN(\RegFile/_1349_ ) );
AOI22_X1 \RegFile/_5384_ ( .A1(\RegFile/_1340_ ), .A2(\RegFile/_1349_ ), .B1(\RegFile/_0104_ ), .B2(\RegFile/_1198_ ), .ZN(\RegFile/_0669_ ) );
NAND3_X1 \RegFile/_5385_ ( .A1(\RegFile/_0761_ ), .A2(\RegFile/_3433_ ), .A3(\RegFile/_0765_ ), .ZN(\RegFile/_1350_ ) );
NAND3_X1 \RegFile/_5386_ ( .A1(\RegFile/_0801_ ), .A2(\RegFile/_0784_ ), .A3(\RegFile/_3689_ ), .ZN(\RegFile/_1351_ ) );
AND2_X1 \RegFile/_5387_ ( .A1(\RegFile/_1350_ ), .A2(\RegFile/_1351_ ), .ZN(\RegFile/_1352_ ) );
INV_X1 \RegFile/_5388_ ( .A(\RegFile/_3657_ ), .ZN(\RegFile/_1353_ ) );
OAI221_X1 \RegFile/_5389_ ( .A(\RegFile/_1352_ ), .B1(\RegFile/_0791_ ), .B2(\RegFile/_0107_ ), .C1(\RegFile/_1353_ ), .C2(\RegFile/_0901_ ), .ZN(\RegFile/_1354_ ) );
AND3_X1 \RegFile/_5390_ ( .A1(\RegFile/_0961_ ), .A2(\RegFile/_3369_ ), .A3(\RegFile/_0834_ ), .ZN(\RegFile/_1355_ ) );
NAND3_X1 \RegFile/_5391_ ( .A1(\RegFile/_0841_ ), .A2(\RegFile/_3529_ ), .A3(\RegFile/_0787_ ), .ZN(\RegFile/_1356_ ) );
NAND3_X1 \RegFile/_5392_ ( .A1(\RegFile/_0842_ ), .A2(\RegFile/_0836_ ), .A3(\RegFile/_3401_ ), .ZN(\RegFile/_1357_ ) );
NAND2_X1 \RegFile/_5393_ ( .A1(\RegFile/_1356_ ), .A2(\RegFile/_1357_ ), .ZN(\RegFile/_1358_ ) );
AND3_X1 \RegFile/_5394_ ( .A1(\RegFile/_0844_ ), .A2(\RegFile/_0784_ ), .A3(\RegFile/_3337_ ), .ZN(\RegFile/_1359_ ) );
NOR4_X1 \RegFile/_5395_ ( .A1(\RegFile/_1354_ ), .A2(\RegFile/_1355_ ), .A3(\RegFile/_1358_ ), .A4(\RegFile/_1359_ ), .ZN(\RegFile/_1360_ ) );
NAND3_X1 \RegFile/_5396_ ( .A1(\RegFile/_0825_ ), .A2(\RegFile/_3753_ ), .A3(\RegFile/_0770_ ), .ZN(\RegFile/_1361_ ) );
AND3_X1 \RegFile/_5397_ ( .A1(\RegFile/_0800_ ), .A2(\RegFile/_3625_ ), .A3(\RegFile/_0768_ ), .ZN(\RegFile/_1362_ ) );
AOI221_X4 \RegFile/_5398_ ( .A(\RegFile/_1362_ ), .B1(\RegFile/_3593_ ), .B2(\RegFile/_0779_ ), .C1(\RegFile/_3561_ ), .C2(\RegFile/_0820_ ), .ZN(\RegFile/_1363_ ) );
NAND3_X1 \RegFile/_5399_ ( .A1(\RegFile/_0893_ ), .A2(\RegFile/_3721_ ), .A3(\RegFile/_0894_ ), .ZN(\RegFile/_1364_ ) );
AOI21_X1 \RegFile/_5400_ ( .A(\RegFile/_0807_ ), .B1(\RegFile/_0828_ ), .B2(\RegFile/_3785_ ), .ZN(\RegFile/_1365_ ) );
AND4_X1 \RegFile/_5401_ ( .A1(\RegFile/_1361_ ), .A2(\RegFile/_1363_ ), .A3(\RegFile/_1364_ ), .A4(\RegFile/_1365_ ), .ZN(\RegFile/_1366_ ) );
AOI22_X1 \RegFile/_5402_ ( .A1(\RegFile/_1360_ ), .A2(\RegFile/_1366_ ), .B1(\RegFile/_0106_ ), .B2(\RegFile/_0811_ ), .ZN(\RegFile/_0671_ ) );
NAND3_X1 \RegFile/_5403_ ( .A1(\RegFile/_0785_ ), .A2(\RegFile/_3562_ ), .A3(\RegFile/_0787_ ), .ZN(\RegFile/_1367_ ) );
NAND3_X1 \RegFile/_5404_ ( .A1(\RegFile/_0864_ ), .A2(\RegFile/_3754_ ), .A3(\RegFile/_0769_ ), .ZN(\RegFile/_1368_ ) );
NAND3_X1 \RegFile/_5405_ ( .A1(\RegFile/_0864_ ), .A2(\RegFile/_0761_ ), .A3(\RegFile/_3786_ ), .ZN(\RegFile/_1369_ ) );
NAND3_X1 \RegFile/_5406_ ( .A1(\RegFile/_0801_ ), .A2(\RegFile/_3722_ ), .A3(\RegFile/_0775_ ), .ZN(\RegFile/_1370_ ) );
AND4_X1 \RegFile/_5407_ ( .A1(\RegFile/_0813_ ), .A2(\RegFile/_1368_ ), .A3(\RegFile/_1369_ ), .A4(\RegFile/_1370_ ), .ZN(\RegFile/_1371_ ) );
NAND3_X1 \RegFile/_5408_ ( .A1(\RegFile/_0893_ ), .A2(\RegFile/_3626_ ), .A3(\RegFile/_0891_ ), .ZN(\RegFile/_1372_ ) );
NAND3_X1 \RegFile/_5409_ ( .A1(\RegFile/_0943_ ), .A2(\RegFile/_0787_ ), .A3(\RegFile/_3594_ ), .ZN(\RegFile/_1373_ ) );
AND4_X1 \RegFile/_5410_ ( .A1(\RegFile/_1367_ ), .A2(\RegFile/_1371_ ), .A3(\RegFile/_1372_ ), .A4(\RegFile/_1373_ ), .ZN(\RegFile/_1374_ ) );
NAND3_X1 \RegFile/_5411_ ( .A1(\RegFile/_0825_ ), .A2(\RegFile/_3370_ ), .A3(\RegFile/_0943_ ), .ZN(\RegFile/_1375_ ) );
INV_X1 \RegFile/_5412_ ( .A(\RegFile/_0109_ ), .ZN(\RegFile/_1376_ ) );
NAND3_X1 \RegFile/_5413_ ( .A1(\RegFile/_0755_ ), .A2(\RegFile/_1376_ ), .A3(\RegFile/_0764_ ), .ZN(\RegFile/_1377_ ) );
INV_X1 \RegFile/_5414_ ( .A(\RegFile/_3658_ ), .ZN(\RegFile/_1378_ ) );
OAI21_X1 \RegFile/_5415_ ( .A(\RegFile/_1377_ ), .B1(\RegFile/_0901_ ), .B2(\RegFile/_1378_ ), .ZN(\RegFile/_1379_ ) );
AOI221_X4 \RegFile/_5416_ ( .A(\RegFile/_1379_ ), .B1(\RegFile/_3434_ ), .B2(\RegFile/_0888_ ), .C1(\RegFile/_3690_ ), .C2(\RegFile/_0815_ ), .ZN(\RegFile/_1380_ ) );
NAND3_X1 \RegFile/_5417_ ( .A1(\RegFile/_0954_ ), .A2(\RegFile/_0785_ ), .A3(\RegFile/_3338_ ), .ZN(\RegFile/_1381_ ) );
AOI22_X1 \RegFile/_5418_ ( .A1(\RegFile/_0822_ ), .A2(\RegFile/_3530_ ), .B1(\RegFile/_0872_ ), .B2(\RegFile/_3402_ ), .ZN(\RegFile/_1382_ ) );
AND4_X1 \RegFile/_5419_ ( .A1(\RegFile/_1375_ ), .A2(\RegFile/_1380_ ), .A3(\RegFile/_1381_ ), .A4(\RegFile/_1382_ ), .ZN(\RegFile/_1383_ ) );
AOI22_X1 \RegFile/_5420_ ( .A1(\RegFile/_1374_ ), .A2(\RegFile/_1383_ ), .B1(\RegFile/_0108_ ), .B2(\RegFile/_0811_ ), .ZN(\RegFile/_0672_ ) );
INV_X1 \RegFile/_5421_ ( .A(\RegFile/_0646_ ), .ZN(\RegFile/_1384_ ) );
AND2_X1 \RegFile/_5422_ ( .A1(\RegFile/_1384_ ), .A2(\RegFile/_0647_ ), .ZN(\RegFile/_1385_ ) );
BUF_X4 \RegFile/_5423_ ( .A(\RegFile/_1385_ ), .Z(\RegFile/_1386_ ) );
BUF_X4 \RegFile/_5424_ ( .A(\RegFile/_1386_ ), .Z(\RegFile/_1387_ ) );
NOR2_X2 \RegFile/_5425_ ( .A1(\RegFile/_0645_ ), .A2(\RegFile/_0644_ ), .ZN(\RegFile/_1388_ ) );
BUF_X4 \RegFile/_5426_ ( .A(\RegFile/_1388_ ), .Z(\RegFile/_1389_ ) );
NAND3_X1 \RegFile/_5427_ ( .A1(\RegFile/_1387_ ), .A2(\RegFile/_3730_ ), .A3(\RegFile/_1389_ ), .ZN(\RegFile/_1390_ ) );
INV_X1 \RegFile/_5428_ ( .A(\RegFile/_0645_ ), .ZN(\RegFile/_1391_ ) );
AND2_X2 \RegFile/_5429_ ( .A1(\RegFile/_1391_ ), .A2(\RegFile/_0644_ ), .ZN(\RegFile/_1392_ ) );
BUF_X2 \RegFile/_5430_ ( .A(\RegFile/_1392_ ), .Z(\RegFile/_1393_ ) );
NOR2_X1 \RegFile/_5431_ ( .A1(\RegFile/_0646_ ), .A2(\RegFile/_0647_ ), .ZN(\RegFile/_1394_ ) );
BUF_X2 \RegFile/_5432_ ( .A(\RegFile/_1394_ ), .Z(\RegFile/_1395_ ) );
BUF_X4 \RegFile/_5433_ ( .A(\RegFile/_1395_ ), .Z(\RegFile/_1396_ ) );
NAND3_X1 \RegFile/_5434_ ( .A1(\RegFile/_1393_ ), .A2(\RegFile/_3506_ ), .A3(\RegFile/_1396_ ), .ZN(\RegFile/_1397_ ) );
NOR2_X1 \RegFile/_5435_ ( .A1(\RegFile/_1384_ ), .A2(\RegFile/_0647_ ), .ZN(\RegFile/_1398_ ) );
BUF_X4 \RegFile/_5436_ ( .A(\RegFile/_1398_ ), .Z(\RegFile/_1399_ ) );
NAND3_X1 \RegFile/_5437_ ( .A1(\RegFile/_1399_ ), .A2(\RegFile/_3602_ ), .A3(\RegFile/_1389_ ), .ZN(\RegFile/_1400_ ) );
NOR2_X1 \RegFile/_5438_ ( .A1(\RegFile/_1391_ ), .A2(\RegFile/_0644_ ), .ZN(\RegFile/_1401_ ) );
BUF_X4 \RegFile/_5439_ ( .A(\RegFile/_1401_ ), .Z(\RegFile/_1402_ ) );
BUF_X4 \RegFile/_5440_ ( .A(\RegFile/_1402_ ), .Z(\RegFile/_1403_ ) );
NAND3_X1 \RegFile/_5441_ ( .A1(\RegFile/_1399_ ), .A2(\RegFile/_1403_ ), .A3(\RegFile/_3666_ ), .ZN(\RegFile/_1404_ ) );
AND4_X1 \RegFile/_5442_ ( .A1(\RegFile/_1390_ ), .A2(\RegFile/_1397_ ), .A3(\RegFile/_1400_ ), .A4(\RegFile/_1404_ ), .ZN(\RegFile/_1405_ ) );
AND2_X2 \RegFile/_5443_ ( .A1(\RegFile/_0646_ ), .A2(\RegFile/_0647_ ), .ZN(\RegFile/_1406_ ) );
AND2_X2 \RegFile/_5444_ ( .A1(\RegFile/_1401_ ), .A2(\RegFile/_1406_ ), .ZN(\RegFile/_1407_ ) );
INV_X1 \RegFile/_5445_ ( .A(\RegFile/_1407_ ), .ZN(\RegFile/_1408_ ) );
BUF_X4 \RegFile/_5446_ ( .A(\RegFile/_1408_ ), .Z(\RegFile/_1409_ ) );
NOR2_X1 \RegFile/_5447_ ( .A1(\RegFile/_1409_ ), .A2(\RegFile/_0111_ ), .ZN(\RegFile/_1410_ ) );
AND2_X2 \RegFile/_5448_ ( .A1(\RegFile/_1401_ ), .A2(\RegFile/_1394_ ), .ZN(\RegFile/_1411_ ) );
BUF_X4 \RegFile/_5449_ ( .A(\RegFile/_1411_ ), .Z(\RegFile/_1412_ ) );
AOI21_X1 \RegFile/_5450_ ( .A(\RegFile/_1410_ ), .B1(\RegFile/_3538_ ), .B2(\RegFile/_1412_ ), .ZN(\RegFile/_1413_ ) );
AND2_X2 \RegFile/_5451_ ( .A1(\RegFile/_0645_ ), .A2(\RegFile/_0644_ ), .ZN(\RegFile/_1414_ ) );
AND2_X1 \RegFile/_5452_ ( .A1(\RegFile/_1406_ ), .A2(\RegFile/_1414_ ), .ZN(\RegFile/_1415_ ) );
BUF_X4 \RegFile/_5453_ ( .A(\RegFile/_1415_ ), .Z(\RegFile/_1416_ ) );
BUF_X4 \RegFile/_5454_ ( .A(\RegFile/_1416_ ), .Z(\RegFile/_1417_ ) );
INV_X1 \RegFile/_5455_ ( .A(\RegFile/_1417_ ), .ZN(\RegFile/_1418_ ) );
BUF_X2 \RegFile/_5456_ ( .A(\RegFile/_1399_ ), .Z(\RegFile/_1419_ ) );
BUF_X4 \RegFile/_5457_ ( .A(\RegFile/_1419_ ), .Z(\RegFile/_1420_ ) );
BUF_X4 \RegFile/_5458_ ( .A(\RegFile/_1414_ ), .Z(\RegFile/_1421_ ) );
BUF_X4 \RegFile/_5459_ ( .A(\RegFile/_1421_ ), .Z(\RegFile/_1422_ ) );
NAND3_X1 \RegFile/_5460_ ( .A1(\RegFile/_1420_ ), .A2(\RegFile/_3698_ ), .A3(\RegFile/_1422_ ), .ZN(\RegFile/_1423_ ) );
AND4_X1 \RegFile/_5461_ ( .A1(\RegFile/_1405_ ), .A2(\RegFile/_1413_ ), .A3(\RegFile/_1418_ ), .A4(\RegFile/_1423_ ), .ZN(\RegFile/_1424_ ) );
AND3_X1 \RegFile/_5462_ ( .A1(\RegFile/_1385_ ), .A2(\RegFile/_1402_ ), .A3(\RegFile/_3314_ ), .ZN(\RegFile/_1425_ ) );
AND2_X2 \RegFile/_5463_ ( .A1(\RegFile/_1385_ ), .A2(\RegFile/_1392_ ), .ZN(\RegFile/_1426_ ) );
AND2_X2 \RegFile/_5464_ ( .A1(\RegFile/_1392_ ), .A2(\RegFile/_1398_ ), .ZN(\RegFile/_1427_ ) );
AOI221_X4 \RegFile/_5465_ ( .A(\RegFile/_1425_ ), .B1(\RegFile/_1426_ ), .B2(\RegFile/_3762_ ), .C1(\RegFile/_3634_ ), .C2(\RegFile/_1427_ ), .ZN(\RegFile/_1428_ ) );
BUF_X2 \RegFile/_5466_ ( .A(\RegFile/_1392_ ), .Z(\RegFile/_1429_ ) );
BUF_X4 \RegFile/_5467_ ( .A(\RegFile/_1429_ ), .Z(\RegFile/_1430_ ) );
BUF_X4 \RegFile/_5468_ ( .A(\RegFile/_1406_ ), .Z(\RegFile/_1431_ ) );
BUF_X4 \RegFile/_5469_ ( .A(\RegFile/_1431_ ), .Z(\RegFile/_1432_ ) );
NAND3_X1 \RegFile/_5470_ ( .A1(\RegFile/_1430_ ), .A2(\RegFile/_3410_ ), .A3(\RegFile/_1432_ ), .ZN(\RegFile/_1433_ ) );
BUF_X4 \RegFile/_5471_ ( .A(\RegFile/_1389_ ), .Z(\RegFile/_1434_ ) );
NAND3_X1 \RegFile/_5472_ ( .A1(\RegFile/_1432_ ), .A2(\RegFile/_1434_ ), .A3(\RegFile/_3378_ ), .ZN(\RegFile/_1435_ ) );
AND2_X1 \RegFile/_5473_ ( .A1(\RegFile/_1385_ ), .A2(\RegFile/_1414_ ), .ZN(\RegFile/_1436_ ) );
BUF_X4 \RegFile/_5474_ ( .A(\RegFile/_1436_ ), .Z(\RegFile/_1437_ ) );
AND2_X1 \RegFile/_5475_ ( .A1(\RegFile/_1414_ ), .A2(\RegFile/_1394_ ), .ZN(\RegFile/_1438_ ) );
AOI22_X1 \RegFile/_5476_ ( .A1(\RegFile/_1437_ ), .A2(\RegFile/_3346_ ), .B1(\RegFile/_1438_ ), .B2(\RegFile/_3570_ ), .ZN(\RegFile/_1439_ ) );
AND4_X1 \RegFile/_5477_ ( .A1(\RegFile/_1428_ ), .A2(\RegFile/_1433_ ), .A3(\RegFile/_1435_ ), .A4(\RegFile/_1439_ ), .ZN(\RegFile/_1440_ ) );
BUF_X4 \RegFile/_5478_ ( .A(\RegFile/_1416_ ), .Z(\RegFile/_1441_ ) );
BUF_X4 \RegFile/_5479_ ( .A(\RegFile/_1441_ ), .Z(\RegFile/_1442_ ) );
AOI22_X1 \RegFile/_5480_ ( .A1(\RegFile/_1424_ ), .A2(\RegFile/_1440_ ), .B1(\RegFile/_0110_ ), .B2(\RegFile/_1442_ ), .ZN(\RegFile/_0680_ ) );
BUF_X4 \RegFile/_5481_ ( .A(\RegFile/_1386_ ), .Z(\RegFile/_1443_ ) );
AND2_X2 \RegFile/_5482_ ( .A1(\RegFile/_1443_ ), .A2(\RegFile/_1403_ ), .ZN(\RegFile/_1444_ ) );
AOI22_X1 \RegFile/_5483_ ( .A1(\RegFile/_3325_ ), .A2(\RegFile/_1444_ ), .B1(\RegFile/_1437_ ), .B2(\RegFile/_3357_ ), .ZN(\RegFile/_1445_ ) );
NOR2_X1 \RegFile/_5484_ ( .A1(\RegFile/_1409_ ), .A2(\RegFile/_0113_ ), .ZN(\RegFile/_1446_ ) );
AND2_X2 \RegFile/_5485_ ( .A1(\RegFile/_1399_ ), .A2(\RegFile/_1388_ ), .ZN(\RegFile/_1447_ ) );
BUF_X4 \RegFile/_5486_ ( .A(\RegFile/_1447_ ), .Z(\RegFile/_1448_ ) );
AOI21_X1 \RegFile/_5487_ ( .A(\RegFile/_1446_ ), .B1(\RegFile/_3613_ ), .B2(\RegFile/_1448_ ), .ZN(\RegFile/_1449_ ) );
AND2_X2 \RegFile/_5488_ ( .A1(\RegFile/_1392_ ), .A2(\RegFile/_1395_ ), .ZN(\RegFile/_1450_ ) );
AND2_X1 \RegFile/_5489_ ( .A1(\RegFile/_1406_ ), .A2(\RegFile/_1388_ ), .ZN(\RegFile/_1451_ ) );
AOI22_X1 \RegFile/_5490_ ( .A1(\RegFile/_1450_ ), .A2(\RegFile/_3517_ ), .B1(\RegFile/_1451_ ), .B2(\RegFile/_3389_ ), .ZN(\RegFile/_1452_ ) );
AOI22_X1 \RegFile/_5491_ ( .A1(\RegFile/_1412_ ), .A2(\RegFile/_3549_ ), .B1(\RegFile/_1438_ ), .B2(\RegFile/_3581_ ), .ZN(\RegFile/_1453_ ) );
AND4_X1 \RegFile/_5492_ ( .A1(\RegFile/_1445_ ), .A2(\RegFile/_1449_ ), .A3(\RegFile/_1452_ ), .A4(\RegFile/_1453_ ), .ZN(\RegFile/_1454_ ) );
BUF_X2 \RegFile/_5493_ ( .A(\RegFile/_1393_ ), .Z(\RegFile/_1455_ ) );
NAND3_X1 \RegFile/_5494_ ( .A1(\RegFile/_1455_ ), .A2(\RegFile/_1419_ ), .A3(\RegFile/_3645_ ), .ZN(\RegFile/_1456_ ) );
AND2_X1 \RegFile/_5495_ ( .A1(\RegFile/_1398_ ), .A2(\RegFile/_1401_ ), .ZN(\RegFile/_1457_ ) );
INV_X1 \RegFile/_5496_ ( .A(\RegFile/_1457_ ), .ZN(\RegFile/_1458_ ) );
INV_X1 \RegFile/_5497_ ( .A(\RegFile/_3421_ ), .ZN(\RegFile/_1459_ ) );
AND2_X2 \RegFile/_5498_ ( .A1(\RegFile/_1392_ ), .A2(\RegFile/_1406_ ), .ZN(\RegFile/_1460_ ) );
BUF_X4 \RegFile/_5499_ ( .A(\RegFile/_1460_ ), .Z(\RegFile/_1461_ ) );
INV_X1 \RegFile/_5500_ ( .A(\RegFile/_1461_ ), .ZN(\RegFile/_1462_ ) );
OAI221_X1 \RegFile/_5501_ ( .A(\RegFile/_1456_ ), .B1(\RegFile/_1458_ ), .B2(\RegFile/_0817_ ), .C1(\RegFile/_1459_ ), .C2(\RegFile/_1462_ ), .ZN(\RegFile/_1463_ ) );
BUF_X4 \RegFile/_5502_ ( .A(\RegFile/_1388_ ), .Z(\RegFile/_1464_ ) );
NAND4_X1 \RegFile/_5503_ ( .A1(\RegFile/_1464_ ), .A2(\RegFile/_3741_ ), .A3(\RegFile/_1384_ ), .A4(\RegFile/_0647_ ), .ZN(\RegFile/_1465_ ) );
NAND2_X2 \RegFile/_5504_ ( .A1(\RegFile/_1399_ ), .A2(\RegFile/_1421_ ), .ZN(\RegFile/_1466_ ) );
OAI21_X1 \RegFile/_5505_ ( .A(\RegFile/_1465_ ), .B1(\RegFile/_1466_ ), .B2(\RegFile/_0849_ ), .ZN(\RegFile/_1467_ ) );
BUF_X2 \RegFile/_5506_ ( .A(\RegFile/_1386_ ), .Z(\RegFile/_1468_ ) );
AND3_X1 \RegFile/_5507_ ( .A1(\RegFile/_1468_ ), .A2(\RegFile/_1429_ ), .A3(\RegFile/_3773_ ), .ZN(\RegFile/_1469_ ) );
NOR4_X1 \RegFile/_5508_ ( .A1(\RegFile/_1463_ ), .A2(\RegFile/_1441_ ), .A3(\RegFile/_1467_ ), .A4(\RegFile/_1469_ ), .ZN(\RegFile/_1470_ ) );
AOI22_X1 \RegFile/_5509_ ( .A1(\RegFile/_1454_ ), .A2(\RegFile/_1470_ ), .B1(\RegFile/_0112_ ), .B2(\RegFile/_1442_ ), .ZN(\RegFile/_0691_ ) );
BUF_X4 \RegFile/_5510_ ( .A(\RegFile/_1403_ ), .Z(\RegFile/_1471_ ) );
BUF_X4 \RegFile/_5511_ ( .A(\RegFile/_1396_ ), .Z(\RegFile/_1472_ ) );
NAND3_X1 \RegFile/_5512_ ( .A1(\RegFile/_1471_ ), .A2(\RegFile/_3560_ ), .A3(\RegFile/_1472_ ), .ZN(\RegFile/_1473_ ) );
INV_X1 \RegFile/_5513_ ( .A(\RegFile/_1438_ ), .ZN(\RegFile/_1474_ ) );
INV_X1 \RegFile/_5514_ ( .A(\RegFile/_3592_ ), .ZN(\RegFile/_1475_ ) );
INV_X1 \RegFile/_5515_ ( .A(\RegFile/_1448_ ), .ZN(\RegFile/_1476_ ) );
BUF_X4 \RegFile/_5516_ ( .A(\RegFile/_1476_ ), .Z(\RegFile/_1477_ ) );
INV_X1 \RegFile/_5517_ ( .A(\RegFile/_3624_ ), .ZN(\RegFile/_1478_ ) );
OAI221_X1 \RegFile/_5518_ ( .A(\RegFile/_1473_ ), .B1(\RegFile/_1474_ ), .B2(\RegFile/_1475_ ), .C1(\RegFile/_1477_ ), .C2(\RegFile/_1478_ ), .ZN(\RegFile/_1479_ ) );
BUF_X4 \RegFile/_5519_ ( .A(\RegFile/_1417_ ), .Z(\RegFile/_1480_ ) );
CLKBUF_X2 \RegFile/_5520_ ( .A(\RegFile/_1386_ ), .Z(\RegFile/_1481_ ) );
CLKBUF_X2 \RegFile/_5521_ ( .A(\RegFile/_1393_ ), .Z(\RegFile/_1482_ ) );
AND3_X1 \RegFile/_5522_ ( .A1(\RegFile/_1481_ ), .A2(\RegFile/_1482_ ), .A3(\RegFile/_3784_ ), .ZN(\RegFile/_1483_ ) );
BUF_X2 \RegFile/_5523_ ( .A(\RegFile/_1388_ ), .Z(\RegFile/_1484_ ) );
NAND3_X1 \RegFile/_5524_ ( .A1(\RegFile/_1468_ ), .A2(\RegFile/_3752_ ), .A3(\RegFile/_1484_ ), .ZN(\RegFile/_1485_ ) );
BUF_X4 \RegFile/_5525_ ( .A(\RegFile/_1466_ ), .Z(\RegFile/_1486_ ) );
OAI21_X1 \RegFile/_5526_ ( .A(\RegFile/_1485_ ), .B1(\RegFile/_1486_ ), .B2(\RegFile/_0859_ ), .ZN(\RegFile/_1487_ ) );
NOR4_X1 \RegFile/_5527_ ( .A1(\RegFile/_1479_ ), .A2(\RegFile/_1480_ ), .A3(\RegFile/_1483_ ), .A4(\RegFile/_1487_ ), .ZN(\RegFile/_1488_ ) );
BUF_X4 \RegFile/_5528_ ( .A(\RegFile/_1403_ ), .Z(\RegFile/_1489_ ) );
NAND3_X1 \RegFile/_5529_ ( .A1(\RegFile/_1420_ ), .A2(\RegFile/_1489_ ), .A3(\RegFile/_3688_ ), .ZN(\RegFile/_1490_ ) );
NAND3_X1 \RegFile/_5530_ ( .A1(\RegFile/_1393_ ), .A2(\RegFile/_3528_ ), .A3(\RegFile/_1396_ ), .ZN(\RegFile/_1491_ ) );
NAND3_X1 \RegFile/_5531_ ( .A1(\RegFile/_1443_ ), .A2(\RegFile/_1403_ ), .A3(\RegFile/_3336_ ), .ZN(\RegFile/_1492_ ) );
NAND3_X1 \RegFile/_5532_ ( .A1(\RegFile/_1443_ ), .A2(\RegFile/_3368_ ), .A3(\RegFile/_1421_ ), .ZN(\RegFile/_1493_ ) );
NAND3_X1 \RegFile/_5533_ ( .A1(\RegFile/_1431_ ), .A2(\RegFile/_1389_ ), .A3(\RegFile/_3400_ ), .ZN(\RegFile/_1494_ ) );
AND4_X1 \RegFile/_5534_ ( .A1(\RegFile/_1491_ ), .A2(\RegFile/_1492_ ), .A3(\RegFile/_1493_ ), .A4(\RegFile/_1494_ ), .ZN(\RegFile/_1495_ ) );
NAND3_X1 \RegFile/_5535_ ( .A1(\RegFile/_1430_ ), .A2(\RegFile/_3432_ ), .A3(\RegFile/_1432_ ), .ZN(\RegFile/_1496_ ) );
AOI22_X1 \RegFile/_5536_ ( .A1(\RegFile/_3656_ ), .A2(\RegFile/_1427_ ), .B1(\RegFile/_1407_ ), .B2(\RegFile/_0867_ ), .ZN(\RegFile/_1497_ ) );
AND4_X1 \RegFile/_5537_ ( .A1(\RegFile/_1490_ ), .A2(\RegFile/_1495_ ), .A3(\RegFile/_1496_ ), .A4(\RegFile/_1497_ ), .ZN(\RegFile/_1498_ ) );
AOI22_X1 \RegFile/_5538_ ( .A1(\RegFile/_1488_ ), .A2(\RegFile/_1498_ ), .B1(\RegFile/_0114_ ), .B2(\RegFile/_1442_ ), .ZN(\RegFile/_0702_ ) );
NAND3_X1 \RegFile/_5539_ ( .A1(\RegFile/_1430_ ), .A2(\RegFile/_3531_ ), .A3(\RegFile/_1472_ ), .ZN(\RegFile/_1499_ ) );
INV_X1 \RegFile/_5540_ ( .A(\RegFile/_1427_ ), .ZN(\RegFile/_1500_ ) );
INV_X1 \RegFile/_5541_ ( .A(\RegFile/_3659_ ), .ZN(\RegFile/_1501_ ) );
OAI22_X1 \RegFile/_5542_ ( .A1(\RegFile/_1500_ ), .A2(\RegFile/_1501_ ), .B1(\RegFile/_1408_ ), .B2(\RegFile/_0117_ ), .ZN(\RegFile/_1502_ ) );
AOI221_X4 \RegFile/_5543_ ( .A(\RegFile/_1502_ ), .B1(\RegFile/_3435_ ), .B2(\RegFile/_1460_ ), .C1(\RegFile/_3691_ ), .C2(\RegFile/_1457_ ), .ZN(\RegFile/_1503_ ) );
NAND3_X1 \RegFile/_5544_ ( .A1(\RegFile/_1432_ ), .A2(\RegFile/_1434_ ), .A3(\RegFile/_3403_ ), .ZN(\RegFile/_1504_ ) );
AOI22_X1 \RegFile/_5545_ ( .A1(\RegFile/_3339_ ), .A2(\RegFile/_1444_ ), .B1(\RegFile/_1437_ ), .B2(\RegFile/_3371_ ), .ZN(\RegFile/_1505_ ) );
AND4_X1 \RegFile/_5546_ ( .A1(\RegFile/_1499_ ), .A2(\RegFile/_1503_ ), .A3(\RegFile/_1504_ ), .A4(\RegFile/_1505_ ), .ZN(\RegFile/_1506_ ) );
BUF_X4 \RegFile/_5547_ ( .A(\RegFile/_1421_ ), .Z(\RegFile/_1507_ ) );
CLKBUF_X2 \RegFile/_5548_ ( .A(\RegFile/_1396_ ), .Z(\RegFile/_1508_ ) );
NAND3_X1 \RegFile/_5549_ ( .A1(\RegFile/_1507_ ), .A2(\RegFile/_1508_ ), .A3(\RegFile/_3595_ ), .ZN(\RegFile/_1509_ ) );
INV_X1 \RegFile/_5550_ ( .A(\RegFile/_3627_ ), .ZN(\RegFile/_1510_ ) );
INV_X1 \RegFile/_5551_ ( .A(\RegFile/_3563_ ), .ZN(\RegFile/_1511_ ) );
INV_X2 \RegFile/_5552_ ( .A(\RegFile/_1412_ ), .ZN(\RegFile/_1512_ ) );
OAI221_X1 \RegFile/_5553_ ( .A(\RegFile/_1509_ ), .B1(\RegFile/_1477_ ), .B2(\RegFile/_1510_ ), .C1(\RegFile/_1511_ ), .C2(\RegFile/_1512_ ), .ZN(\RegFile/_1513_ ) );
NAND3_X1 \RegFile/_5554_ ( .A1(\RegFile/_1387_ ), .A2(\RegFile/_3755_ ), .A3(\RegFile/_1464_ ), .ZN(\RegFile/_1514_ ) );
INV_X1 \RegFile/_5555_ ( .A(\RegFile/_3723_ ), .ZN(\RegFile/_1515_ ) );
OAI21_X1 \RegFile/_5556_ ( .A(\RegFile/_1514_ ), .B1(\RegFile/_1466_ ), .B2(\RegFile/_1515_ ), .ZN(\RegFile/_1516_ ) );
AND3_X1 \RegFile/_5557_ ( .A1(\RegFile/_1468_ ), .A2(\RegFile/_1429_ ), .A3(\RegFile/_3787_ ), .ZN(\RegFile/_1517_ ) );
NOR4_X1 \RegFile/_5558_ ( .A1(\RegFile/_1513_ ), .A2(\RegFile/_1441_ ), .A3(\RegFile/_1516_ ), .A4(\RegFile/_1517_ ), .ZN(\RegFile/_1518_ ) );
AOI22_X1 \RegFile/_5559_ ( .A1(\RegFile/_1506_ ), .A2(\RegFile/_1518_ ), .B1(\RegFile/_0116_ ), .B2(\RegFile/_1442_ ), .ZN(\RegFile/_0705_ ) );
BUF_X4 \RegFile/_5560_ ( .A(\RegFile/_1457_ ), .Z(\RegFile/_1519_ ) );
AOI22_X1 \RegFile/_5561_ ( .A1(\RegFile/_3692_ ), .A2(\RegFile/_1519_ ), .B1(\RegFile/_1461_ ), .B2(\RegFile/_3436_ ), .ZN(\RegFile/_1520_ ) );
BUF_X4 \RegFile/_5562_ ( .A(\RegFile/_1409_ ), .Z(\RegFile/_1521_ ) );
BUF_X4 \RegFile/_5563_ ( .A(\RegFile/_1500_ ), .Z(\RegFile/_1522_ ) );
OAI221_X1 \RegFile/_5564_ ( .A(\RegFile/_1520_ ), .B1(\RegFile/_1521_ ), .B2(\RegFile/_0119_ ), .C1(\RegFile/_0902_ ), .C2(\RegFile/_1522_ ), .ZN(\RegFile/_1523_ ) );
BUF_X2 \RegFile/_5565_ ( .A(\RegFile/_1393_ ), .Z(\RegFile/_1524_ ) );
AND3_X1 \RegFile/_5566_ ( .A1(\RegFile/_1524_ ), .A2(\RegFile/_3532_ ), .A3(\RegFile/_1508_ ), .ZN(\RegFile/_1525_ ) );
BUF_X2 \RegFile/_5567_ ( .A(\RegFile/_1431_ ), .Z(\RegFile/_1526_ ) );
CLKBUF_X2 \RegFile/_5568_ ( .A(\RegFile/_1388_ ), .Z(\RegFile/_1527_ ) );
AND3_X1 \RegFile/_5569_ ( .A1(\RegFile/_1526_ ), .A2(\RegFile/_3404_ ), .A3(\RegFile/_1527_ ), .ZN(\RegFile/_1528_ ) );
BUF_X4 \RegFile/_5570_ ( .A(\RegFile/_1443_ ), .Z(\RegFile/_1529_ ) );
BUF_X4 \RegFile/_5571_ ( .A(\RegFile/_1403_ ), .Z(\RegFile/_1530_ ) );
NAND3_X1 \RegFile/_5572_ ( .A1(\RegFile/_1529_ ), .A2(\RegFile/_1530_ ), .A3(\RegFile/_3340_ ), .ZN(\RegFile/_1531_ ) );
BUF_X2 \RegFile/_5573_ ( .A(\RegFile/_1421_ ), .Z(\RegFile/_1532_ ) );
NAND3_X1 \RegFile/_5574_ ( .A1(\RegFile/_1481_ ), .A2(\RegFile/_3372_ ), .A3(\RegFile/_1532_ ), .ZN(\RegFile/_1533_ ) );
NAND2_X1 \RegFile/_5575_ ( .A1(\RegFile/_1531_ ), .A2(\RegFile/_1533_ ), .ZN(\RegFile/_1534_ ) );
NOR4_X1 \RegFile/_5576_ ( .A1(\RegFile/_1523_ ), .A2(\RegFile/_1525_ ), .A3(\RegFile/_1528_ ), .A4(\RegFile/_1534_ ), .ZN(\RegFile/_1535_ ) );
BUF_X2 \RegFile/_5577_ ( .A(\RegFile/_1395_ ), .Z(\RegFile/_1536_ ) );
NAND3_X1 \RegFile/_5578_ ( .A1(\RegFile/_1532_ ), .A2(\RegFile/_1536_ ), .A3(\RegFile/_3596_ ), .ZN(\RegFile/_1537_ ) );
OAI221_X1 \RegFile/_5579_ ( .A(\RegFile/_1537_ ), .B1(\RegFile/_1476_ ), .B2(\RegFile/_0910_ ), .C1(\RegFile/_0915_ ), .C2(\RegFile/_1512_ ), .ZN(\RegFile/_1538_ ) );
CLKBUF_X2 \RegFile/_5580_ ( .A(\RegFile/_1386_ ), .Z(\RegFile/_1539_ ) );
AND3_X1 \RegFile/_5581_ ( .A1(\RegFile/_1539_ ), .A2(\RegFile/_1429_ ), .A3(\RegFile/_3788_ ), .ZN(\RegFile/_1540_ ) );
NAND3_X1 \RegFile/_5582_ ( .A1(\RegFile/_1387_ ), .A2(\RegFile/_3756_ ), .A3(\RegFile/_1389_ ), .ZN(\RegFile/_1541_ ) );
OAI21_X1 \RegFile/_5583_ ( .A(\RegFile/_1541_ ), .B1(\RegFile/_1466_ ), .B2(\RegFile/_0905_ ), .ZN(\RegFile/_1542_ ) );
NOR4_X1 \RegFile/_5584_ ( .A1(\RegFile/_1538_ ), .A2(\RegFile/_1441_ ), .A3(\RegFile/_1540_ ), .A4(\RegFile/_1542_ ), .ZN(\RegFile/_1543_ ) );
AOI22_X1 \RegFile/_5585_ ( .A1(\RegFile/_1535_ ), .A2(\RegFile/_1543_ ), .B1(\RegFile/_0118_ ), .B2(\RegFile/_1442_ ), .ZN(\RegFile/_0706_ ) );
NAND3_X1 \RegFile/_5586_ ( .A1(\RegFile/_1507_ ), .A2(\RegFile/_1472_ ), .A3(\RegFile/_3597_ ), .ZN(\RegFile/_1544_ ) );
INV_X1 \RegFile/_5587_ ( .A(\RegFile/_3629_ ), .ZN(\RegFile/_1545_ ) );
INV_X1 \RegFile/_5588_ ( .A(\RegFile/_3565_ ), .ZN(\RegFile/_1546_ ) );
OAI221_X1 \RegFile/_5589_ ( .A(\RegFile/_1544_ ), .B1(\RegFile/_1477_ ), .B2(\RegFile/_1545_ ), .C1(\RegFile/_1546_ ), .C2(\RegFile/_1512_ ), .ZN(\RegFile/_1547_ ) );
NAND3_X1 \RegFile/_5590_ ( .A1(\RegFile/_1539_ ), .A2(\RegFile/_3757_ ), .A3(\RegFile/_1484_ ), .ZN(\RegFile/_1548_ ) );
INV_X1 \RegFile/_5591_ ( .A(\RegFile/_3725_ ), .ZN(\RegFile/_1549_ ) );
OAI21_X1 \RegFile/_5592_ ( .A(\RegFile/_1548_ ), .B1(\RegFile/_1486_ ), .B2(\RegFile/_1549_ ), .ZN(\RegFile/_1550_ ) );
AND3_X1 \RegFile/_5593_ ( .A1(\RegFile/_1539_ ), .A2(\RegFile/_1482_ ), .A3(\RegFile/_3789_ ), .ZN(\RegFile/_1551_ ) );
NOR4_X1 \RegFile/_5594_ ( .A1(\RegFile/_1547_ ), .A2(\RegFile/_1480_ ), .A3(\RegFile/_1550_ ), .A4(\RegFile/_1551_ ), .ZN(\RegFile/_1552_ ) );
INV_X1 \RegFile/_5595_ ( .A(\RegFile/_3661_ ), .ZN(\RegFile/_1553_ ) );
OAI22_X1 \RegFile/_5596_ ( .A1(\RegFile/_1522_ ), .A2(\RegFile/_1553_ ), .B1(\RegFile/_1521_ ), .B2(\RegFile/_0121_ ), .ZN(\RegFile/_1554_ ) );
BUF_X4 \RegFile/_5597_ ( .A(\RegFile/_1386_ ), .Z(\RegFile/_1555_ ) );
BUF_X2 \RegFile/_5598_ ( .A(\RegFile/_1402_ ), .Z(\RegFile/_1556_ ) );
NAND3_X1 \RegFile/_5599_ ( .A1(\RegFile/_1555_ ), .A2(\RegFile/_1556_ ), .A3(\RegFile/_3341_ ), .ZN(\RegFile/_1557_ ) );
CLKBUF_X2 \RegFile/_5600_ ( .A(\RegFile/_1392_ ), .Z(\RegFile/_1558_ ) );
NAND3_X1 \RegFile/_5601_ ( .A1(\RegFile/_1558_ ), .A2(\RegFile/_3533_ ), .A3(\RegFile/_1536_ ), .ZN(\RegFile/_1559_ ) );
BUF_X4 \RegFile/_5602_ ( .A(\RegFile/_1421_ ), .Z(\RegFile/_1560_ ) );
NAND3_X1 \RegFile/_5603_ ( .A1(\RegFile/_1387_ ), .A2(\RegFile/_3373_ ), .A3(\RegFile/_1560_ ), .ZN(\RegFile/_1561_ ) );
CLKBUF_X2 \RegFile/_5604_ ( .A(\RegFile/_1406_ ), .Z(\RegFile/_1562_ ) );
NAND3_X1 \RegFile/_5605_ ( .A1(\RegFile/_1562_ ), .A2(\RegFile/_1464_ ), .A3(\RegFile/_3405_ ), .ZN(\RegFile/_1563_ ) );
NAND4_X1 \RegFile/_5606_ ( .A1(\RegFile/_1557_ ), .A2(\RegFile/_1559_ ), .A3(\RegFile/_1561_ ), .A4(\RegFile/_1563_ ), .ZN(\RegFile/_1564_ ) );
AND3_X1 \RegFile/_5607_ ( .A1(\RegFile/_1419_ ), .A2(\RegFile/_1556_ ), .A3(\RegFile/_3693_ ), .ZN(\RegFile/_1565_ ) );
AND3_X1 \RegFile/_5608_ ( .A1(\RegFile/_1558_ ), .A2(\RegFile/_3437_ ), .A3(\RegFile/_1562_ ), .ZN(\RegFile/_1566_ ) );
NOR4_X1 \RegFile/_5609_ ( .A1(\RegFile/_1554_ ), .A2(\RegFile/_1564_ ), .A3(\RegFile/_1565_ ), .A4(\RegFile/_1566_ ), .ZN(\RegFile/_1567_ ) );
AOI22_X1 \RegFile/_5610_ ( .A1(\RegFile/_1552_ ), .A2(\RegFile/_1567_ ), .B1(\RegFile/_0120_ ), .B2(\RegFile/_1442_ ), .ZN(\RegFile/_0707_ ) );
NAND3_X1 \RegFile/_5611_ ( .A1(\RegFile/_1471_ ), .A2(\RegFile/_3566_ ), .A3(\RegFile/_1472_ ), .ZN(\RegFile/_1568_ ) );
INV_X1 \RegFile/_5612_ ( .A(\RegFile/_3598_ ), .ZN(\RegFile/_1569_ ) );
INV_X1 \RegFile/_5613_ ( .A(\RegFile/_3630_ ), .ZN(\RegFile/_1570_ ) );
OAI221_X1 \RegFile/_5614_ ( .A(\RegFile/_1568_ ), .B1(\RegFile/_1474_ ), .B2(\RegFile/_1569_ ), .C1(\RegFile/_1477_ ), .C2(\RegFile/_1570_ ), .ZN(\RegFile/_1571_ ) );
AND3_X1 \RegFile/_5615_ ( .A1(\RegFile/_1481_ ), .A2(\RegFile/_1482_ ), .A3(\RegFile/_3790_ ), .ZN(\RegFile/_1572_ ) );
NAND3_X1 \RegFile/_5616_ ( .A1(\RegFile/_1468_ ), .A2(\RegFile/_3758_ ), .A3(\RegFile/_1484_ ), .ZN(\RegFile/_1573_ ) );
INV_X1 \RegFile/_5617_ ( .A(\RegFile/_3726_ ), .ZN(\RegFile/_1574_ ) );
OAI21_X1 \RegFile/_5618_ ( .A(\RegFile/_1573_ ), .B1(\RegFile/_1486_ ), .B2(\RegFile/_1574_ ), .ZN(\RegFile/_1575_ ) );
NOR4_X1 \RegFile/_5619_ ( .A1(\RegFile/_1571_ ), .A2(\RegFile/_1480_ ), .A3(\RegFile/_1572_ ), .A4(\RegFile/_1575_ ), .ZN(\RegFile/_1576_ ) );
BUF_X4 \RegFile/_5620_ ( .A(\RegFile/_1399_ ), .Z(\RegFile/_1577_ ) );
NAND3_X1 \RegFile/_5621_ ( .A1(\RegFile/_1524_ ), .A2(\RegFile/_1577_ ), .A3(\RegFile/_3662_ ), .ZN(\RegFile/_1578_ ) );
NAND3_X1 \RegFile/_5622_ ( .A1(\RegFile/_1455_ ), .A2(\RegFile/_3438_ ), .A3(\RegFile/_1526_ ), .ZN(\RegFile/_1579_ ) );
NAND3_X1 \RegFile/_5623_ ( .A1(\RegFile/_1471_ ), .A2(\RegFile/_0951_ ), .A3(\RegFile/_1526_ ), .ZN(\RegFile/_1580_ ) );
NAND3_X1 \RegFile/_5624_ ( .A1(\RegFile/_1419_ ), .A2(\RegFile/_1530_ ), .A3(\RegFile/_3694_ ), .ZN(\RegFile/_1581_ ) );
NAND4_X1 \RegFile/_5625_ ( .A1(\RegFile/_1578_ ), .A2(\RegFile/_1579_ ), .A3(\RegFile/_1580_ ), .A4(\RegFile/_1581_ ), .ZN(\RegFile/_1582_ ) );
BUF_X2 \RegFile/_5626_ ( .A(\RegFile/_1386_ ), .Z(\RegFile/_1583_ ) );
NAND3_X1 \RegFile/_5627_ ( .A1(\RegFile/_1583_ ), .A2(\RegFile/_1471_ ), .A3(\RegFile/_3342_ ), .ZN(\RegFile/_1584_ ) );
NAND3_X1 \RegFile/_5628_ ( .A1(\RegFile/_1529_ ), .A2(\RegFile/_3374_ ), .A3(\RegFile/_1532_ ), .ZN(\RegFile/_1585_ ) );
NAND2_X1 \RegFile/_5629_ ( .A1(\RegFile/_1584_ ), .A2(\RegFile/_1585_ ), .ZN(\RegFile/_1586_ ) );
AND3_X1 \RegFile/_5630_ ( .A1(\RegFile/_1482_ ), .A2(\RegFile/_3534_ ), .A3(\RegFile/_1536_ ), .ZN(\RegFile/_1587_ ) );
CLKBUF_X2 \RegFile/_5631_ ( .A(\RegFile/_1431_ ), .Z(\RegFile/_1588_ ) );
AND3_X1 \RegFile/_5632_ ( .A1(\RegFile/_1588_ ), .A2(\RegFile/_3406_ ), .A3(\RegFile/_1484_ ), .ZN(\RegFile/_1589_ ) );
NOR4_X1 \RegFile/_5633_ ( .A1(\RegFile/_1582_ ), .A2(\RegFile/_1586_ ), .A3(\RegFile/_1587_ ), .A4(\RegFile/_1589_ ), .ZN(\RegFile/_1590_ ) );
AOI22_X1 \RegFile/_5634_ ( .A1(\RegFile/_1576_ ), .A2(\RegFile/_1590_ ), .B1(\RegFile/_0122_ ), .B2(\RegFile/_1442_ ), .ZN(\RegFile/_0708_ ) );
NAND3_X1 \RegFile/_5635_ ( .A1(\RegFile/_1399_ ), .A2(\RegFile/_1402_ ), .A3(\RegFile/_3695_ ), .ZN(\RegFile/_1591_ ) );
OAI21_X1 \RegFile/_5636_ ( .A(\RegFile/_1591_ ), .B1(\RegFile/_1409_ ), .B2(\RegFile/_0125_ ), .ZN(\RegFile/_1592_ ) );
AOI221_X4 \RegFile/_5637_ ( .A(\RegFile/_1592_ ), .B1(\RegFile/_3567_ ), .B2(\RegFile/_1411_ ), .C1(\RegFile/_3535_ ), .C2(\RegFile/_1450_ ), .ZN(\RegFile/_1593_ ) );
BUF_X4 \RegFile/_5638_ ( .A(\RegFile/_1426_ ), .Z(\RegFile/_1594_ ) );
AOI21_X1 \RegFile/_5639_ ( .A(\RegFile/_1416_ ), .B1(\RegFile/_1594_ ), .B2(\RegFile/_3791_ ), .ZN(\RegFile/_1595_ ) );
BUF_X4 \RegFile/_5640_ ( .A(\RegFile/_1387_ ), .Z(\RegFile/_1596_ ) );
NAND3_X1 \RegFile/_5641_ ( .A1(\RegFile/_1596_ ), .A2(\RegFile/_3759_ ), .A3(\RegFile/_1434_ ), .ZN(\RegFile/_1597_ ) );
NAND3_X1 \RegFile/_5642_ ( .A1(\RegFile/_1430_ ), .A2(\RegFile/_1420_ ), .A3(\RegFile/_3663_ ), .ZN(\RegFile/_1598_ ) );
AND4_X1 \RegFile/_5643_ ( .A1(\RegFile/_1593_ ), .A2(\RegFile/_1595_ ), .A3(\RegFile/_1597_ ), .A4(\RegFile/_1598_ ), .ZN(\RegFile/_1599_ ) );
CLKBUF_X2 \RegFile/_5644_ ( .A(\RegFile/_1414_ ), .Z(\RegFile/_1600_ ) );
AND3_X1 \RegFile/_5645_ ( .A1(\RegFile/_1600_ ), .A2(\RegFile/_3599_ ), .A3(\RegFile/_1395_ ), .ZN(\RegFile/_1601_ ) );
AOI221_X4 \RegFile/_5646_ ( .A(\RegFile/_1601_ ), .B1(\RegFile/_1448_ ), .B2(\RegFile/_3631_ ), .C1(\RegFile/_3375_ ), .C2(\RegFile/_1437_ ), .ZN(\RegFile/_1602_ ) );
AND3_X1 \RegFile/_5647_ ( .A1(\RegFile/_1393_ ), .A2(\RegFile/_3439_ ), .A3(\RegFile/_1431_ ), .ZN(\RegFile/_1603_ ) );
AOI21_X1 \RegFile/_5648_ ( .A(\RegFile/_1603_ ), .B1(\RegFile/_3343_ ), .B2(\RegFile/_1444_ ), .ZN(\RegFile/_1604_ ) );
NAND3_X1 \RegFile/_5649_ ( .A1(\RegFile/_1432_ ), .A2(\RegFile/_1434_ ), .A3(\RegFile/_3407_ ), .ZN(\RegFile/_1605_ ) );
BUF_X4 \RegFile/_5650_ ( .A(\RegFile/_1399_ ), .Z(\RegFile/_1606_ ) );
NAND3_X1 \RegFile/_5651_ ( .A1(\RegFile/_1606_ ), .A2(\RegFile/_3727_ ), .A3(\RegFile/_1422_ ), .ZN(\RegFile/_1607_ ) );
AND4_X1 \RegFile/_5652_ ( .A1(\RegFile/_1602_ ), .A2(\RegFile/_1604_ ), .A3(\RegFile/_1605_ ), .A4(\RegFile/_1607_ ), .ZN(\RegFile/_1608_ ) );
AOI22_X1 \RegFile/_5653_ ( .A1(\RegFile/_1599_ ), .A2(\RegFile/_1608_ ), .B1(\RegFile/_0124_ ), .B2(\RegFile/_1442_ ), .ZN(\RegFile/_0709_ ) );
AOI22_X1 \RegFile/_5654_ ( .A1(\RegFile/_3696_ ), .A2(\RegFile/_1519_ ), .B1(\RegFile/_1461_ ), .B2(\RegFile/_3440_ ), .ZN(\RegFile/_1609_ ) );
OAI221_X1 \RegFile/_5655_ ( .A(\RegFile/_1609_ ), .B1(\RegFile/_1521_ ), .B2(\RegFile/_0127_ ), .C1(\RegFile/_0977_ ), .C2(\RegFile/_1522_ ), .ZN(\RegFile/_1610_ ) );
AND3_X1 \RegFile/_5656_ ( .A1(\RegFile/_1524_ ), .A2(\RegFile/_3536_ ), .A3(\RegFile/_1508_ ), .ZN(\RegFile/_1611_ ) );
AND3_X1 \RegFile/_5657_ ( .A1(\RegFile/_1588_ ), .A2(\RegFile/_3408_ ), .A3(\RegFile/_1527_ ), .ZN(\RegFile/_1612_ ) );
NAND3_X1 \RegFile/_5658_ ( .A1(\RegFile/_1529_ ), .A2(\RegFile/_1530_ ), .A3(\RegFile/_3344_ ), .ZN(\RegFile/_1613_ ) );
NAND3_X1 \RegFile/_5659_ ( .A1(\RegFile/_1481_ ), .A2(\RegFile/_3376_ ), .A3(\RegFile/_1532_ ), .ZN(\RegFile/_1614_ ) );
NAND2_X1 \RegFile/_5660_ ( .A1(\RegFile/_1613_ ), .A2(\RegFile/_1614_ ), .ZN(\RegFile/_1615_ ) );
NOR4_X1 \RegFile/_5661_ ( .A1(\RegFile/_1610_ ), .A2(\RegFile/_1611_ ), .A3(\RegFile/_1612_ ), .A4(\RegFile/_1615_ ), .ZN(\RegFile/_1616_ ) );
AOI21_X1 \RegFile/_5662_ ( .A(\RegFile/_1417_ ), .B1(\RegFile/_1594_ ), .B2(\RegFile/_3792_ ), .ZN(\RegFile/_1617_ ) );
AND3_X1 \RegFile/_5663_ ( .A1(\RegFile/_1600_ ), .A2(\RegFile/_3600_ ), .A3(\RegFile/_1394_ ), .ZN(\RegFile/_1618_ ) );
AOI221_X4 \RegFile/_5664_ ( .A(\RegFile/_1618_ ), .B1(\RegFile/_1447_ ), .B2(\RegFile/_3632_ ), .C1(\RegFile/_3568_ ), .C2(\RegFile/_1412_ ), .ZN(\RegFile/_1619_ ) );
BUF_X4 \RegFile/_5665_ ( .A(\RegFile/_1389_ ), .Z(\RegFile/_1620_ ) );
NAND3_X1 \RegFile/_5666_ ( .A1(\RegFile/_1583_ ), .A2(\RegFile/_3760_ ), .A3(\RegFile/_1620_ ), .ZN(\RegFile/_1621_ ) );
NAND3_X1 \RegFile/_5667_ ( .A1(\RegFile/_1606_ ), .A2(\RegFile/_3728_ ), .A3(\RegFile/_1422_ ), .ZN(\RegFile/_1622_ ) );
AND4_X1 \RegFile/_5668_ ( .A1(\RegFile/_1617_ ), .A2(\RegFile/_1619_ ), .A3(\RegFile/_1621_ ), .A4(\RegFile/_1622_ ), .ZN(\RegFile/_1623_ ) );
AOI22_X1 \RegFile/_5669_ ( .A1(\RegFile/_1616_ ), .A2(\RegFile/_1623_ ), .B1(\RegFile/_0126_ ), .B2(\RegFile/_1442_ ), .ZN(\RegFile/_0710_ ) );
NOR2_X1 \RegFile/_5670_ ( .A1(\RegFile/_1409_ ), .A2(\RegFile/_0065_ ), .ZN(\RegFile/_1624_ ) );
AOI221_X4 \RegFile/_5671_ ( .A(\RegFile/_1624_ ), .B1(\RegFile/_3377_ ), .B2(\RegFile/_1437_ ), .C1(\RegFile/_3665_ ), .C2(\RegFile/_1427_ ), .ZN(\RegFile/_1625_ ) );
NAND3_X1 \RegFile/_5672_ ( .A1(\RegFile/_1596_ ), .A2(\RegFile/_1489_ ), .A3(\RegFile/_3345_ ), .ZN(\RegFile/_1626_ ) );
NAND3_X1 \RegFile/_5673_ ( .A1(\RegFile/_1489_ ), .A2(\RegFile/_3569_ ), .A3(\RegFile/_1472_ ), .ZN(\RegFile/_1627_ ) );
AOI22_X1 \RegFile/_5674_ ( .A1(\RegFile/_1426_ ), .A2(\RegFile/_3793_ ), .B1(\RegFile/_1451_ ), .B2(\RegFile/_3409_ ), .ZN(\RegFile/_1628_ ) );
AND4_X1 \RegFile/_5675_ ( .A1(\RegFile/_1625_ ), .A2(\RegFile/_1626_ ), .A3(\RegFile/_1627_ ), .A4(\RegFile/_1628_ ), .ZN(\RegFile/_1629_ ) );
AOI22_X1 \RegFile/_5676_ ( .A1(\RegFile/_1450_ ), .A2(\RegFile/_3537_ ), .B1(\RegFile/_1457_ ), .B2(\RegFile/_3697_ ), .ZN(\RegFile/_1630_ ) );
NAND3_X1 \RegFile/_5677_ ( .A1(\RegFile/_1532_ ), .A2(\RegFile/_1536_ ), .A3(\RegFile/_3601_ ), .ZN(\RegFile/_1631_ ) );
OAI211_X2 \RegFile/_5678_ ( .A(\RegFile/_1630_ ), .B(\RegFile/_1631_ ), .C1(\RegFile/_1004_ ), .C2(\RegFile/_1477_ ), .ZN(\RegFile/_1632_ ) );
NAND4_X1 \RegFile/_5679_ ( .A1(\RegFile/_1389_ ), .A2(\RegFile/_3761_ ), .A3(\RegFile/_1384_ ), .A4(\RegFile/_0647_ ), .ZN(\RegFile/_1633_ ) );
OAI21_X1 \RegFile/_5680_ ( .A(\RegFile/_1633_ ), .B1(\RegFile/_1466_ ), .B2(\RegFile/_1009_ ), .ZN(\RegFile/_1634_ ) );
AND3_X1 \RegFile/_5681_ ( .A1(\RegFile/_1558_ ), .A2(\RegFile/_3441_ ), .A3(\RegFile/_1562_ ), .ZN(\RegFile/_1635_ ) );
NOR4_X1 \RegFile/_5682_ ( .A1(\RegFile/_1632_ ), .A2(\RegFile/_1441_ ), .A3(\RegFile/_1634_ ), .A4(\RegFile/_1635_ ), .ZN(\RegFile/_1636_ ) );
AOI22_X1 \RegFile/_5683_ ( .A1(\RegFile/_1629_ ), .A2(\RegFile/_1636_ ), .B1(\RegFile/_0064_ ), .B2(\RegFile/_1442_ ), .ZN(\RegFile/_0711_ ) );
AOI22_X1 \RegFile/_5684_ ( .A1(\RegFile/_3667_ ), .A2(\RegFile/_1519_ ), .B1(\RegFile/_1461_ ), .B2(\RegFile/_3411_ ), .ZN(\RegFile/_1637_ ) );
OAI221_X1 \RegFile/_5685_ ( .A(\RegFile/_1637_ ), .B1(\RegFile/_1521_ ), .B2(\RegFile/_0067_ ), .C1(\RegFile/_1014_ ), .C2(\RegFile/_1522_ ), .ZN(\RegFile/_1638_ ) );
AND3_X1 \RegFile/_5686_ ( .A1(\RegFile/_1524_ ), .A2(\RegFile/_3507_ ), .A3(\RegFile/_1508_ ), .ZN(\RegFile/_1639_ ) );
AND3_X1 \RegFile/_5687_ ( .A1(\RegFile/_1588_ ), .A2(\RegFile/_3379_ ), .A3(\RegFile/_1527_ ), .ZN(\RegFile/_1640_ ) );
NAND3_X1 \RegFile/_5688_ ( .A1(\RegFile/_1529_ ), .A2(\RegFile/_1530_ ), .A3(\RegFile/_3315_ ), .ZN(\RegFile/_1641_ ) );
NAND3_X1 \RegFile/_5689_ ( .A1(\RegFile/_1555_ ), .A2(\RegFile/_3347_ ), .A3(\RegFile/_1560_ ), .ZN(\RegFile/_1642_ ) );
NAND2_X1 \RegFile/_5690_ ( .A1(\RegFile/_1641_ ), .A2(\RegFile/_1642_ ), .ZN(\RegFile/_1643_ ) );
NOR4_X1 \RegFile/_5691_ ( .A1(\RegFile/_1638_ ), .A2(\RegFile/_1639_ ), .A3(\RegFile/_1640_ ), .A4(\RegFile/_1643_ ), .ZN(\RegFile/_1644_ ) );
AOI21_X1 \RegFile/_5692_ ( .A(\RegFile/_1417_ ), .B1(\RegFile/_1594_ ), .B2(\RegFile/_3763_ ), .ZN(\RegFile/_1645_ ) );
AND3_X1 \RegFile/_5693_ ( .A1(\RegFile/_1600_ ), .A2(\RegFile/_3571_ ), .A3(\RegFile/_1394_ ), .ZN(\RegFile/_1646_ ) );
AOI221_X4 \RegFile/_5694_ ( .A(\RegFile/_1646_ ), .B1(\RegFile/_1447_ ), .B2(\RegFile/_3603_ ), .C1(\RegFile/_3539_ ), .C2(\RegFile/_1411_ ), .ZN(\RegFile/_1647_ ) );
NAND3_X1 \RegFile/_5695_ ( .A1(\RegFile/_1583_ ), .A2(\RegFile/_3731_ ), .A3(\RegFile/_1620_ ), .ZN(\RegFile/_1648_ ) );
NAND3_X1 \RegFile/_5696_ ( .A1(\RegFile/_1606_ ), .A2(\RegFile/_3699_ ), .A3(\RegFile/_1422_ ), .ZN(\RegFile/_1649_ ) );
AND4_X1 \RegFile/_5697_ ( .A1(\RegFile/_1645_ ), .A2(\RegFile/_1647_ ), .A3(\RegFile/_1648_ ), .A4(\RegFile/_1649_ ), .ZN(\RegFile/_1650_ ) );
BUF_X4 \RegFile/_5698_ ( .A(\RegFile/_1441_ ), .Z(\RegFile/_1651_ ) );
AOI22_X1 \RegFile/_5699_ ( .A1(\RegFile/_1644_ ), .A2(\RegFile/_1650_ ), .B1(\RegFile/_0066_ ), .B2(\RegFile/_1651_ ), .ZN(\RegFile/_0681_ ) );
NAND3_X1 \RegFile/_5700_ ( .A1(\RegFile/_1507_ ), .A2(\RegFile/_1472_ ), .A3(\RegFile/_3572_ ), .ZN(\RegFile/_1652_ ) );
INV_X1 \RegFile/_5701_ ( .A(\RegFile/_3604_ ), .ZN(\RegFile/_1653_ ) );
INV_X1 \RegFile/_5702_ ( .A(\RegFile/_3540_ ), .ZN(\RegFile/_1654_ ) );
OAI221_X1 \RegFile/_5703_ ( .A(\RegFile/_1652_ ), .B1(\RegFile/_1477_ ), .B2(\RegFile/_1653_ ), .C1(\RegFile/_1654_ ), .C2(\RegFile/_1512_ ), .ZN(\RegFile/_1655_ ) );
NAND3_X1 \RegFile/_5704_ ( .A1(\RegFile/_1539_ ), .A2(\RegFile/_3732_ ), .A3(\RegFile/_1484_ ), .ZN(\RegFile/_1656_ ) );
INV_X1 \RegFile/_5705_ ( .A(\RegFile/_3700_ ), .ZN(\RegFile/_1657_ ) );
OAI21_X1 \RegFile/_5706_ ( .A(\RegFile/_1656_ ), .B1(\RegFile/_1486_ ), .B2(\RegFile/_1657_ ), .ZN(\RegFile/_1658_ ) );
AND3_X1 \RegFile/_5707_ ( .A1(\RegFile/_1539_ ), .A2(\RegFile/_1558_ ), .A3(\RegFile/_3764_ ), .ZN(\RegFile/_1659_ ) );
NOR4_X1 \RegFile/_5708_ ( .A1(\RegFile/_1655_ ), .A2(\RegFile/_1480_ ), .A3(\RegFile/_1658_ ), .A4(\RegFile/_1659_ ), .ZN(\RegFile/_1660_ ) );
INV_X1 \RegFile/_5709_ ( .A(\RegFile/_3636_ ), .ZN(\RegFile/_1661_ ) );
OAI22_X1 \RegFile/_5710_ ( .A1(\RegFile/_1522_ ), .A2(\RegFile/_1661_ ), .B1(\RegFile/_1521_ ), .B2(\RegFile/_0069_ ), .ZN(\RegFile/_1662_ ) );
NAND3_X1 \RegFile/_5711_ ( .A1(\RegFile/_1555_ ), .A2(\RegFile/_1556_ ), .A3(\RegFile/_3316_ ), .ZN(\RegFile/_1663_ ) );
NAND3_X1 \RegFile/_5712_ ( .A1(\RegFile/_1429_ ), .A2(\RegFile/_3508_ ), .A3(\RegFile/_1536_ ), .ZN(\RegFile/_1664_ ) );
NAND3_X1 \RegFile/_5713_ ( .A1(\RegFile/_1387_ ), .A2(\RegFile/_3348_ ), .A3(\RegFile/_1560_ ), .ZN(\RegFile/_1665_ ) );
NAND3_X1 \RegFile/_5714_ ( .A1(\RegFile/_1562_ ), .A2(\RegFile/_1464_ ), .A3(\RegFile/_3380_ ), .ZN(\RegFile/_1666_ ) );
NAND4_X1 \RegFile/_5715_ ( .A1(\RegFile/_1663_ ), .A2(\RegFile/_1664_ ), .A3(\RegFile/_1665_ ), .A4(\RegFile/_1666_ ), .ZN(\RegFile/_1667_ ) );
AND3_X1 \RegFile/_5716_ ( .A1(\RegFile/_1419_ ), .A2(\RegFile/_1556_ ), .A3(\RegFile/_3668_ ), .ZN(\RegFile/_1668_ ) );
AND3_X1 \RegFile/_5717_ ( .A1(\RegFile/_1558_ ), .A2(\RegFile/_3412_ ), .A3(\RegFile/_1562_ ), .ZN(\RegFile/_1669_ ) );
NOR4_X1 \RegFile/_5718_ ( .A1(\RegFile/_1662_ ), .A2(\RegFile/_1667_ ), .A3(\RegFile/_1668_ ), .A4(\RegFile/_1669_ ), .ZN(\RegFile/_1670_ ) );
AOI22_X1 \RegFile/_5719_ ( .A1(\RegFile/_1660_ ), .A2(\RegFile/_1670_ ), .B1(\RegFile/_0068_ ), .B2(\RegFile/_1651_ ), .ZN(\RegFile/_0682_ ) );
AOI22_X1 \RegFile/_5720_ ( .A1(\RegFile/_3669_ ), .A2(\RegFile/_1519_ ), .B1(\RegFile/_1461_ ), .B2(\RegFile/_3413_ ), .ZN(\RegFile/_1671_ ) );
OAI221_X1 \RegFile/_5721_ ( .A(\RegFile/_1671_ ), .B1(\RegFile/_1521_ ), .B2(\RegFile/_0071_ ), .C1(\RegFile/_1049_ ), .C2(\RegFile/_1522_ ), .ZN(\RegFile/_1672_ ) );
AND3_X1 \RegFile/_5722_ ( .A1(\RegFile/_1455_ ), .A2(\RegFile/_3509_ ), .A3(\RegFile/_1508_ ), .ZN(\RegFile/_1673_ ) );
AND3_X1 \RegFile/_5723_ ( .A1(\RegFile/_1588_ ), .A2(\RegFile/_3381_ ), .A3(\RegFile/_1527_ ), .ZN(\RegFile/_1674_ ) );
NAND3_X1 \RegFile/_5724_ ( .A1(\RegFile/_1529_ ), .A2(\RegFile/_1530_ ), .A3(\RegFile/_3317_ ), .ZN(\RegFile/_1675_ ) );
NAND3_X1 \RegFile/_5725_ ( .A1(\RegFile/_1555_ ), .A2(\RegFile/_3349_ ), .A3(\RegFile/_1560_ ), .ZN(\RegFile/_1676_ ) );
NAND2_X1 \RegFile/_5726_ ( .A1(\RegFile/_1675_ ), .A2(\RegFile/_1676_ ), .ZN(\RegFile/_1677_ ) );
NOR4_X1 \RegFile/_5727_ ( .A1(\RegFile/_1672_ ), .A2(\RegFile/_1673_ ), .A3(\RegFile/_1674_ ), .A4(\RegFile/_1677_ ), .ZN(\RegFile/_1678_ ) );
NAND3_X1 \RegFile/_5728_ ( .A1(\RegFile/_1532_ ), .A2(\RegFile/_1536_ ), .A3(\RegFile/_3573_ ), .ZN(\RegFile/_1679_ ) );
OAI221_X1 \RegFile/_5729_ ( .A(\RegFile/_1679_ ), .B1(\RegFile/_1476_ ), .B2(\RegFile/_1056_ ), .C1(\RegFile/_1059_ ), .C2(\RegFile/_1512_ ), .ZN(\RegFile/_1680_ ) );
AND3_X1 \RegFile/_5730_ ( .A1(\RegFile/_1539_ ), .A2(\RegFile/_1429_ ), .A3(\RegFile/_3765_ ), .ZN(\RegFile/_1681_ ) );
NAND3_X1 \RegFile/_5731_ ( .A1(\RegFile/_1387_ ), .A2(\RegFile/_3733_ ), .A3(\RegFile/_1389_ ), .ZN(\RegFile/_1682_ ) );
OAI21_X1 \RegFile/_5732_ ( .A(\RegFile/_1682_ ), .B1(\RegFile/_1466_ ), .B2(\RegFile/_1052_ ), .ZN(\RegFile/_1683_ ) );
NOR4_X1 \RegFile/_5733_ ( .A1(\RegFile/_1680_ ), .A2(\RegFile/_1441_ ), .A3(\RegFile/_1681_ ), .A4(\RegFile/_1683_ ), .ZN(\RegFile/_1684_ ) );
AOI22_X1 \RegFile/_5734_ ( .A1(\RegFile/_1678_ ), .A2(\RegFile/_1684_ ), .B1(\RegFile/_0070_ ), .B2(\RegFile/_1651_ ), .ZN(\RegFile/_0683_ ) );
NAND3_X1 \RegFile/_5735_ ( .A1(\RegFile/_1399_ ), .A2(\RegFile/_1402_ ), .A3(\RegFile/_3670_ ), .ZN(\RegFile/_1685_ ) );
OAI21_X1 \RegFile/_5736_ ( .A(\RegFile/_1685_ ), .B1(\RegFile/_1409_ ), .B2(\RegFile/_0073_ ), .ZN(\RegFile/_1686_ ) );
AOI221_X4 \RegFile/_5737_ ( .A(\RegFile/_1686_ ), .B1(\RegFile/_3766_ ), .B2(\RegFile/_1426_ ), .C1(\RegFile/_3510_ ), .C2(\RegFile/_1450_ ), .ZN(\RegFile/_1687_ ) );
NAND3_X1 \RegFile/_5738_ ( .A1(\RegFile/_1596_ ), .A2(\RegFile/_3734_ ), .A3(\RegFile/_1434_ ), .ZN(\RegFile/_1688_ ) );
AOI22_X1 \RegFile/_5739_ ( .A1(\RegFile/_3606_ ), .A2(\RegFile/_1448_ ), .B1(\RegFile/_1412_ ), .B2(\RegFile/_3542_ ), .ZN(\RegFile/_1689_ ) );
AND4_X1 \RegFile/_5740_ ( .A1(\RegFile/_1418_ ), .A2(\RegFile/_1687_ ), .A3(\RegFile/_1688_ ), .A4(\RegFile/_1689_ ), .ZN(\RegFile/_1690_ ) );
NAND3_X1 \RegFile/_5741_ ( .A1(\RegFile/_1596_ ), .A2(\RegFile/_3350_ ), .A3(\RegFile/_1422_ ), .ZN(\RegFile/_1691_ ) );
NAND3_X1 \RegFile/_5742_ ( .A1(\RegFile/_1385_ ), .A2(\RegFile/_1402_ ), .A3(\RegFile/_3318_ ), .ZN(\RegFile/_1692_ ) );
NAND3_X1 \RegFile/_5743_ ( .A1(\RegFile/_1392_ ), .A2(\RegFile/_3414_ ), .A3(\RegFile/_1406_ ), .ZN(\RegFile/_1693_ ) );
NAND2_X1 \RegFile/_5744_ ( .A1(\RegFile/_1692_ ), .A2(\RegFile/_1693_ ), .ZN(\RegFile/_1694_ ) );
AOI221_X4 \RegFile/_5745_ ( .A(\RegFile/_1694_ ), .B1(\RegFile/_3382_ ), .B2(\RegFile/_1451_ ), .C1(\RegFile/_3574_ ), .C2(\RegFile/_1438_ ), .ZN(\RegFile/_1695_ ) );
NAND3_X1 \RegFile/_5746_ ( .A1(\RegFile/_1420_ ), .A2(\RegFile/_3702_ ), .A3(\RegFile/_1422_ ), .ZN(\RegFile/_1696_ ) );
NAND3_X1 \RegFile/_5747_ ( .A1(\RegFile/_1430_ ), .A2(\RegFile/_1577_ ), .A3(\RegFile/_3638_ ), .ZN(\RegFile/_1697_ ) );
AND4_X1 \RegFile/_5748_ ( .A1(\RegFile/_1691_ ), .A2(\RegFile/_1695_ ), .A3(\RegFile/_1696_ ), .A4(\RegFile/_1697_ ), .ZN(\RegFile/_1698_ ) );
AOI22_X1 \RegFile/_5749_ ( .A1(\RegFile/_1690_ ), .A2(\RegFile/_1698_ ), .B1(\RegFile/_0072_ ), .B2(\RegFile/_1651_ ), .ZN(\RegFile/_0684_ ) );
NAND3_X1 \RegFile/_5750_ ( .A1(\RegFile/_1507_ ), .A2(\RegFile/_1472_ ), .A3(\RegFile/_3575_ ), .ZN(\RegFile/_1699_ ) );
INV_X1 \RegFile/_5751_ ( .A(\RegFile/_3607_ ), .ZN(\RegFile/_1700_ ) );
INV_X1 \RegFile/_5752_ ( .A(\RegFile/_3543_ ), .ZN(\RegFile/_1701_ ) );
OAI221_X1 \RegFile/_5753_ ( .A(\RegFile/_1699_ ), .B1(\RegFile/_1477_ ), .B2(\RegFile/_1700_ ), .C1(\RegFile/_1701_ ), .C2(\RegFile/_1512_ ), .ZN(\RegFile/_1702_ ) );
AND3_X1 \RegFile/_5754_ ( .A1(\RegFile/_1481_ ), .A2(\RegFile/_1482_ ), .A3(\RegFile/_3767_ ), .ZN(\RegFile/_1703_ ) );
NAND3_X1 \RegFile/_5755_ ( .A1(\RegFile/_1468_ ), .A2(\RegFile/_3735_ ), .A3(\RegFile/_1464_ ), .ZN(\RegFile/_1704_ ) );
INV_X1 \RegFile/_5756_ ( .A(\RegFile/_3703_ ), .ZN(\RegFile/_1705_ ) );
OAI21_X1 \RegFile/_5757_ ( .A(\RegFile/_1704_ ), .B1(\RegFile/_1486_ ), .B2(\RegFile/_1705_ ), .ZN(\RegFile/_1706_ ) );
NOR4_X1 \RegFile/_5758_ ( .A1(\RegFile/_1702_ ), .A2(\RegFile/_1480_ ), .A3(\RegFile/_1703_ ), .A4(\RegFile/_1706_ ), .ZN(\RegFile/_1707_ ) );
INV_X1 \RegFile/_5759_ ( .A(\RegFile/_3639_ ), .ZN(\RegFile/_1708_ ) );
OAI22_X1 \RegFile/_5760_ ( .A1(\RegFile/_1522_ ), .A2(\RegFile/_1708_ ), .B1(\RegFile/_1521_ ), .B2(\RegFile/_0075_ ), .ZN(\RegFile/_1709_ ) );
NAND3_X1 \RegFile/_5761_ ( .A1(\RegFile/_1555_ ), .A2(\RegFile/_1556_ ), .A3(\RegFile/_3319_ ), .ZN(\RegFile/_1710_ ) );
NAND3_X1 \RegFile/_5762_ ( .A1(\RegFile/_1429_ ), .A2(\RegFile/_3511_ ), .A3(\RegFile/_1396_ ), .ZN(\RegFile/_1711_ ) );
NAND3_X1 \RegFile/_5763_ ( .A1(\RegFile/_1387_ ), .A2(\RegFile/_3351_ ), .A3(\RegFile/_1560_ ), .ZN(\RegFile/_1712_ ) );
NAND3_X1 \RegFile/_5764_ ( .A1(\RegFile/_1562_ ), .A2(\RegFile/_1464_ ), .A3(\RegFile/_3383_ ), .ZN(\RegFile/_1713_ ) );
NAND4_X1 \RegFile/_5765_ ( .A1(\RegFile/_1710_ ), .A2(\RegFile/_1711_ ), .A3(\RegFile/_1712_ ), .A4(\RegFile/_1713_ ), .ZN(\RegFile/_1714_ ) );
AND3_X1 \RegFile/_5766_ ( .A1(\RegFile/_1419_ ), .A2(\RegFile/_1556_ ), .A3(\RegFile/_3671_ ), .ZN(\RegFile/_1715_ ) );
AND3_X1 \RegFile/_5767_ ( .A1(\RegFile/_1558_ ), .A2(\RegFile/_3415_ ), .A3(\RegFile/_1562_ ), .ZN(\RegFile/_1716_ ) );
NOR4_X1 \RegFile/_5768_ ( .A1(\RegFile/_1709_ ), .A2(\RegFile/_1714_ ), .A3(\RegFile/_1715_ ), .A4(\RegFile/_1716_ ), .ZN(\RegFile/_1717_ ) );
AOI22_X1 \RegFile/_5769_ ( .A1(\RegFile/_1707_ ), .A2(\RegFile/_1717_ ), .B1(\RegFile/_0074_ ), .B2(\RegFile/_1651_ ), .ZN(\RegFile/_0685_ ) );
AND3_X1 \RegFile/_5770_ ( .A1(\RegFile/_1392_ ), .A2(\RegFile/_3512_ ), .A3(\RegFile/_1395_ ), .ZN(\RegFile/_1718_ ) );
NAND3_X1 \RegFile/_5771_ ( .A1(\RegFile/_1402_ ), .A2(\RegFile/_1099_ ), .A3(\RegFile/_1406_ ), .ZN(\RegFile/_1719_ ) );
INV_X1 \RegFile/_5772_ ( .A(\RegFile/_3672_ ), .ZN(\RegFile/_1720_ ) );
OAI21_X1 \RegFile/_5773_ ( .A(\RegFile/_1719_ ), .B1(\RegFile/_1458_ ), .B2(\RegFile/_1720_ ), .ZN(\RegFile/_1721_ ) );
AOI211_X4 \RegFile/_5774_ ( .A(\RegFile/_1718_ ), .B(\RegFile/_1721_ ), .C1(\RegFile/_3544_ ), .C2(\RegFile/_1412_ ), .ZN(\RegFile/_1722_ ) );
AOI21_X1 \RegFile/_5775_ ( .A(\RegFile/_1416_ ), .B1(\RegFile/_1594_ ), .B2(\RegFile/_3768_ ), .ZN(\RegFile/_1723_ ) );
NAND3_X1 \RegFile/_5776_ ( .A1(\RegFile/_1596_ ), .A2(\RegFile/_3736_ ), .A3(\RegFile/_1434_ ), .ZN(\RegFile/_1724_ ) );
NAND3_X1 \RegFile/_5777_ ( .A1(\RegFile/_1430_ ), .A2(\RegFile/_1420_ ), .A3(\RegFile/_3640_ ), .ZN(\RegFile/_1725_ ) );
AND4_X1 \RegFile/_5778_ ( .A1(\RegFile/_1722_ ), .A2(\RegFile/_1723_ ), .A3(\RegFile/_1724_ ), .A4(\RegFile/_1725_ ), .ZN(\RegFile/_1726_ ) );
AND3_X1 \RegFile/_5779_ ( .A1(\RegFile/_1600_ ), .A2(\RegFile/_3576_ ), .A3(\RegFile/_1395_ ), .ZN(\RegFile/_1727_ ) );
AOI221_X4 \RegFile/_5780_ ( .A(\RegFile/_1727_ ), .B1(\RegFile/_1448_ ), .B2(\RegFile/_3608_ ), .C1(\RegFile/_3352_ ), .C2(\RegFile/_1437_ ), .ZN(\RegFile/_1728_ ) );
AOI22_X1 \RegFile/_5781_ ( .A1(\RegFile/_3320_ ), .A2(\RegFile/_1444_ ), .B1(\RegFile/_1461_ ), .B2(\RegFile/_3416_ ), .ZN(\RegFile/_1729_ ) );
NAND3_X1 \RegFile/_5782_ ( .A1(\RegFile/_1432_ ), .A2(\RegFile/_1620_ ), .A3(\RegFile/_3384_ ), .ZN(\RegFile/_1730_ ) );
NAND3_X1 \RegFile/_5783_ ( .A1(\RegFile/_1606_ ), .A2(\RegFile/_3704_ ), .A3(\RegFile/_1422_ ), .ZN(\RegFile/_1731_ ) );
AND4_X1 \RegFile/_5784_ ( .A1(\RegFile/_1728_ ), .A2(\RegFile/_1729_ ), .A3(\RegFile/_1730_ ), .A4(\RegFile/_1731_ ), .ZN(\RegFile/_1732_ ) );
AOI22_X1 \RegFile/_5785_ ( .A1(\RegFile/_1726_ ), .A2(\RegFile/_1732_ ), .B1(\RegFile/_0076_ ), .B2(\RegFile/_1651_ ), .ZN(\RegFile/_0686_ ) );
AOI22_X1 \RegFile/_5786_ ( .A1(\RegFile/_3641_ ), .A2(\RegFile/_1427_ ), .B1(\RegFile/_1407_ ), .B2(\RegFile/_1121_ ), .ZN(\RegFile/_1733_ ) );
INV_X1 \RegFile/_5787_ ( .A(\RegFile/_3417_ ), .ZN(\RegFile/_1734_ ) );
INV_X1 \RegFile/_5788_ ( .A(\RegFile/_3673_ ), .ZN(\RegFile/_1735_ ) );
OAI221_X1 \RegFile/_5789_ ( .A(\RegFile/_1733_ ), .B1(\RegFile/_1462_ ), .B2(\RegFile/_1734_ ), .C1(\RegFile/_1735_ ), .C2(\RegFile/_1458_ ), .ZN(\RegFile/_1736_ ) );
AND3_X1 \RegFile/_5790_ ( .A1(\RegFile/_1455_ ), .A2(\RegFile/_3513_ ), .A3(\RegFile/_1508_ ), .ZN(\RegFile/_1737_ ) );
AND3_X1 \RegFile/_5791_ ( .A1(\RegFile/_1588_ ), .A2(\RegFile/_3385_ ), .A3(\RegFile/_1527_ ), .ZN(\RegFile/_1738_ ) );
NAND3_X1 \RegFile/_5792_ ( .A1(\RegFile/_1529_ ), .A2(\RegFile/_1530_ ), .A3(\RegFile/_3321_ ), .ZN(\RegFile/_1739_ ) );
NAND3_X1 \RegFile/_5793_ ( .A1(\RegFile/_1555_ ), .A2(\RegFile/_3353_ ), .A3(\RegFile/_1560_ ), .ZN(\RegFile/_1740_ ) );
NAND2_X1 \RegFile/_5794_ ( .A1(\RegFile/_1739_ ), .A2(\RegFile/_1740_ ), .ZN(\RegFile/_1741_ ) );
NOR4_X1 \RegFile/_5795_ ( .A1(\RegFile/_1736_ ), .A2(\RegFile/_1737_ ), .A3(\RegFile/_1738_ ), .A4(\RegFile/_1741_ ), .ZN(\RegFile/_1742_ ) );
AOI21_X1 \RegFile/_5796_ ( .A(\RegFile/_1417_ ), .B1(\RegFile/_1594_ ), .B2(\RegFile/_3769_ ), .ZN(\RegFile/_1743_ ) );
AND3_X1 \RegFile/_5797_ ( .A1(\RegFile/_1600_ ), .A2(\RegFile/_3577_ ), .A3(\RegFile/_1394_ ), .ZN(\RegFile/_1744_ ) );
AOI221_X4 \RegFile/_5798_ ( .A(\RegFile/_1744_ ), .B1(\RegFile/_1447_ ), .B2(\RegFile/_3609_ ), .C1(\RegFile/_3545_ ), .C2(\RegFile/_1411_ ), .ZN(\RegFile/_1745_ ) );
NAND3_X1 \RegFile/_5799_ ( .A1(\RegFile/_1583_ ), .A2(\RegFile/_3737_ ), .A3(\RegFile/_1620_ ), .ZN(\RegFile/_1746_ ) );
NAND3_X1 \RegFile/_5800_ ( .A1(\RegFile/_1606_ ), .A2(\RegFile/_3705_ ), .A3(\RegFile/_1422_ ), .ZN(\RegFile/_1747_ ) );
AND4_X1 \RegFile/_5801_ ( .A1(\RegFile/_1743_ ), .A2(\RegFile/_1745_ ), .A3(\RegFile/_1746_ ), .A4(\RegFile/_1747_ ), .ZN(\RegFile/_1748_ ) );
AOI22_X1 \RegFile/_5802_ ( .A1(\RegFile/_1742_ ), .A2(\RegFile/_1748_ ), .B1(\RegFile/_0078_ ), .B2(\RegFile/_1651_ ), .ZN(\RegFile/_0687_ ) );
AOI22_X1 \RegFile/_5803_ ( .A1(\RegFile/_3322_ ), .A2(\RegFile/_1444_ ), .B1(\RegFile/_1437_ ), .B2(\RegFile/_3354_ ), .ZN(\RegFile/_1749_ ) );
NOR2_X1 \RegFile/_5804_ ( .A1(\RegFile/_1409_ ), .A2(\RegFile/_0081_ ), .ZN(\RegFile/_1750_ ) );
AOI21_X1 \RegFile/_5805_ ( .A(\RegFile/_1750_ ), .B1(\RegFile/_3610_ ), .B2(\RegFile/_1448_ ), .ZN(\RegFile/_1751_ ) );
AOI22_X1 \RegFile/_5806_ ( .A1(\RegFile/_1450_ ), .A2(\RegFile/_3514_ ), .B1(\RegFile/_1451_ ), .B2(\RegFile/_3386_ ), .ZN(\RegFile/_1752_ ) );
AOI22_X1 \RegFile/_5807_ ( .A1(\RegFile/_1412_ ), .A2(\RegFile/_3546_ ), .B1(\RegFile/_1438_ ), .B2(\RegFile/_3578_ ), .ZN(\RegFile/_1753_ ) );
AND4_X1 \RegFile/_5808_ ( .A1(\RegFile/_1749_ ), .A2(\RegFile/_1751_ ), .A3(\RegFile/_1752_ ), .A4(\RegFile/_1753_ ), .ZN(\RegFile/_1754_ ) );
NAND3_X1 \RegFile/_5809_ ( .A1(\RegFile/_1524_ ), .A2(\RegFile/_3418_ ), .A3(\RegFile/_1526_ ), .ZN(\RegFile/_1755_ ) );
NAND3_X1 \RegFile/_5810_ ( .A1(\RegFile/_1524_ ), .A2(\RegFile/_1577_ ), .A3(\RegFile/_3642_ ), .ZN(\RegFile/_1756_ ) );
NAND3_X1 \RegFile/_5811_ ( .A1(\RegFile/_1577_ ), .A2(\RegFile/_1489_ ), .A3(\RegFile/_3674_ ), .ZN(\RegFile/_1757_ ) );
NAND3_X1 \RegFile/_5812_ ( .A1(\RegFile/_1755_ ), .A2(\RegFile/_1756_ ), .A3(\RegFile/_1757_ ), .ZN(\RegFile/_1758_ ) );
NAND4_X1 \RegFile/_5813_ ( .A1(\RegFile/_1484_ ), .A2(\RegFile/_3738_ ), .A3(\RegFile/_1384_ ), .A4(\RegFile/_0647_ ), .ZN(\RegFile/_1759_ ) );
OAI21_X1 \RegFile/_5814_ ( .A(\RegFile/_1759_ ), .B1(\RegFile/_1486_ ), .B2(\RegFile/_1141_ ), .ZN(\RegFile/_1760_ ) );
AND3_X1 \RegFile/_5815_ ( .A1(\RegFile/_1539_ ), .A2(\RegFile/_1429_ ), .A3(\RegFile/_3770_ ), .ZN(\RegFile/_1761_ ) );
NOR4_X1 \RegFile/_5816_ ( .A1(\RegFile/_1758_ ), .A2(\RegFile/_1760_ ), .A3(\RegFile/_1761_ ), .A4(\RegFile/_1417_ ), .ZN(\RegFile/_1762_ ) );
AOI22_X1 \RegFile/_5817_ ( .A1(\RegFile/_1754_ ), .A2(\RegFile/_1762_ ), .B1(\RegFile/_0080_ ), .B2(\RegFile/_1651_ ), .ZN(\RegFile/_0688_ ) );
NAND3_X1 \RegFile/_5818_ ( .A1(\RegFile/_1471_ ), .A2(\RegFile/_3547_ ), .A3(\RegFile/_1472_ ), .ZN(\RegFile/_1763_ ) );
INV_X1 \RegFile/_5819_ ( .A(\RegFile/_3579_ ), .ZN(\RegFile/_1764_ ) );
INV_X1 \RegFile/_5820_ ( .A(\RegFile/_3611_ ), .ZN(\RegFile/_1765_ ) );
OAI221_X1 \RegFile/_5821_ ( .A(\RegFile/_1763_ ), .B1(\RegFile/_1474_ ), .B2(\RegFile/_1764_ ), .C1(\RegFile/_1477_ ), .C2(\RegFile/_1765_ ), .ZN(\RegFile/_1766_ ) );
AND3_X1 \RegFile/_5822_ ( .A1(\RegFile/_1481_ ), .A2(\RegFile/_1482_ ), .A3(\RegFile/_3771_ ), .ZN(\RegFile/_1767_ ) );
NAND3_X1 \RegFile/_5823_ ( .A1(\RegFile/_1468_ ), .A2(\RegFile/_3739_ ), .A3(\RegFile/_1464_ ), .ZN(\RegFile/_1768_ ) );
OAI21_X1 \RegFile/_5824_ ( .A(\RegFile/_1768_ ), .B1(\RegFile/_1486_ ), .B2(\RegFile/_1158_ ), .ZN(\RegFile/_1769_ ) );
NOR4_X1 \RegFile/_5825_ ( .A1(\RegFile/_1766_ ), .A2(\RegFile/_1480_ ), .A3(\RegFile/_1767_ ), .A4(\RegFile/_1769_ ), .ZN(\RegFile/_1770_ ) );
NAND3_X1 \RegFile/_5826_ ( .A1(\RegFile/_1524_ ), .A2(\RegFile/_1577_ ), .A3(\RegFile/_3643_ ), .ZN(\RegFile/_1771_ ) );
NAND3_X1 \RegFile/_5827_ ( .A1(\RegFile/_1455_ ), .A2(\RegFile/_3419_ ), .A3(\RegFile/_1526_ ), .ZN(\RegFile/_1772_ ) );
NAND3_X1 \RegFile/_5828_ ( .A1(\RegFile/_1471_ ), .A2(\RegFile/_1149_ ), .A3(\RegFile/_1526_ ), .ZN(\RegFile/_1773_ ) );
NAND3_X1 \RegFile/_5829_ ( .A1(\RegFile/_1419_ ), .A2(\RegFile/_1530_ ), .A3(\RegFile/_3675_ ), .ZN(\RegFile/_1774_ ) );
NAND4_X1 \RegFile/_5830_ ( .A1(\RegFile/_1771_ ), .A2(\RegFile/_1772_ ), .A3(\RegFile/_1773_ ), .A4(\RegFile/_1774_ ), .ZN(\RegFile/_1775_ ) );
NAND3_X1 \RegFile/_5831_ ( .A1(\RegFile/_1583_ ), .A2(\RegFile/_1471_ ), .A3(\RegFile/_3323_ ), .ZN(\RegFile/_1776_ ) );
NAND3_X1 \RegFile/_5832_ ( .A1(\RegFile/_1529_ ), .A2(\RegFile/_3355_ ), .A3(\RegFile/_1532_ ), .ZN(\RegFile/_1777_ ) );
NAND2_X1 \RegFile/_5833_ ( .A1(\RegFile/_1776_ ), .A2(\RegFile/_1777_ ), .ZN(\RegFile/_1778_ ) );
AND3_X1 \RegFile/_5834_ ( .A1(\RegFile/_1482_ ), .A2(\RegFile/_3515_ ), .A3(\RegFile/_1536_ ), .ZN(\RegFile/_1779_ ) );
AND3_X1 \RegFile/_5835_ ( .A1(\RegFile/_1588_ ), .A2(\RegFile/_3387_ ), .A3(\RegFile/_1484_ ), .ZN(\RegFile/_1780_ ) );
NOR4_X1 \RegFile/_5836_ ( .A1(\RegFile/_1775_ ), .A2(\RegFile/_1778_ ), .A3(\RegFile/_1779_ ), .A4(\RegFile/_1780_ ), .ZN(\RegFile/_1781_ ) );
AOI22_X1 \RegFile/_5837_ ( .A1(\RegFile/_1770_ ), .A2(\RegFile/_1781_ ), .B1(\RegFile/_0082_ ), .B2(\RegFile/_1651_ ), .ZN(\RegFile/_0689_ ) );
NAND3_X1 \RegFile/_5838_ ( .A1(\RegFile/_1596_ ), .A2(\RegFile/_3740_ ), .A3(\RegFile/_1434_ ), .ZN(\RegFile/_1782_ ) );
AND3_X1 \RegFile/_5839_ ( .A1(\RegFile/_1600_ ), .A2(\RegFile/_3580_ ), .A3(\RegFile/_1395_ ), .ZN(\RegFile/_1783_ ) );
AOI221_X4 \RegFile/_5840_ ( .A(\RegFile/_1783_ ), .B1(\RegFile/_1448_ ), .B2(\RegFile/_3612_ ), .C1(\RegFile/_3548_ ), .C2(\RegFile/_1412_ ), .ZN(\RegFile/_1784_ ) );
NAND3_X1 \RegFile/_5841_ ( .A1(\RegFile/_1420_ ), .A2(\RegFile/_3708_ ), .A3(\RegFile/_1422_ ), .ZN(\RegFile/_1785_ ) );
AOI21_X1 \RegFile/_5842_ ( .A(\RegFile/_1416_ ), .B1(\RegFile/_1426_ ), .B2(\RegFile/_3772_ ), .ZN(\RegFile/_1786_ ) );
AND4_X1 \RegFile/_5843_ ( .A1(\RegFile/_1782_ ), .A2(\RegFile/_1784_ ), .A3(\RegFile/_1785_ ), .A4(\RegFile/_1786_ ), .ZN(\RegFile/_1787_ ) );
NAND3_X1 \RegFile/_5844_ ( .A1(\RegFile/_1489_ ), .A2(\RegFile/_1162_ ), .A3(\RegFile/_1432_ ), .ZN(\RegFile/_1788_ ) );
AOI22_X1 \RegFile/_5845_ ( .A1(\RegFile/_3676_ ), .A2(\RegFile/_1519_ ), .B1(\RegFile/_1461_ ), .B2(\RegFile/_3420_ ), .ZN(\RegFile/_1789_ ) );
NAND3_X1 \RegFile/_5846_ ( .A1(\RegFile/_1393_ ), .A2(\RegFile/_3516_ ), .A3(\RegFile/_1396_ ), .ZN(\RegFile/_1790_ ) );
NAND3_X1 \RegFile/_5847_ ( .A1(\RegFile/_1443_ ), .A2(\RegFile/_1403_ ), .A3(\RegFile/_3324_ ), .ZN(\RegFile/_1791_ ) );
NAND3_X1 \RegFile/_5848_ ( .A1(\RegFile/_1386_ ), .A2(\RegFile/_3356_ ), .A3(\RegFile/_1421_ ), .ZN(\RegFile/_1792_ ) );
NAND3_X1 \RegFile/_5849_ ( .A1(\RegFile/_1431_ ), .A2(\RegFile/_1388_ ), .A3(\RegFile/_3388_ ), .ZN(\RegFile/_1793_ ) );
AND4_X1 \RegFile/_5850_ ( .A1(\RegFile/_1790_ ), .A2(\RegFile/_1791_ ), .A3(\RegFile/_1792_ ), .A4(\RegFile/_1793_ ), .ZN(\RegFile/_1794_ ) );
NAND3_X1 \RegFile/_5851_ ( .A1(\RegFile/_1524_ ), .A2(\RegFile/_1577_ ), .A3(\RegFile/_3644_ ), .ZN(\RegFile/_1795_ ) );
AND4_X1 \RegFile/_5852_ ( .A1(\RegFile/_1788_ ), .A2(\RegFile/_1789_ ), .A3(\RegFile/_1794_ ), .A4(\RegFile/_1795_ ), .ZN(\RegFile/_1796_ ) );
AOI22_X1 \RegFile/_5853_ ( .A1(\RegFile/_1787_ ), .A2(\RegFile/_1796_ ), .B1(\RegFile/_0084_ ), .B2(\RegFile/_1651_ ), .ZN(\RegFile/_0690_ ) );
AOI22_X1 \RegFile/_5854_ ( .A1(\RegFile/_3646_ ), .A2(\RegFile/_1427_ ), .B1(\RegFile/_1407_ ), .B2(\RegFile/_1193_ ), .ZN(\RegFile/_1797_ ) );
OAI221_X1 \RegFile/_5855_ ( .A(\RegFile/_1797_ ), .B1(\RegFile/_1462_ ), .B2(\RegFile/_1184_ ), .C1(\RegFile/_1183_ ), .C2(\RegFile/_1458_ ), .ZN(\RegFile/_1798_ ) );
AND3_X1 \RegFile/_5856_ ( .A1(\RegFile/_1583_ ), .A2(\RegFile/_3358_ ), .A3(\RegFile/_1532_ ), .ZN(\RegFile/_1799_ ) );
AND3_X1 \RegFile/_5857_ ( .A1(\RegFile/_1481_ ), .A2(\RegFile/_1556_ ), .A3(\RegFile/_3326_ ), .ZN(\RegFile/_1800_ ) );
NAND3_X1 \RegFile/_5858_ ( .A1(\RegFile/_1455_ ), .A2(\RegFile/_3518_ ), .A3(\RegFile/_1536_ ), .ZN(\RegFile/_1801_ ) );
NAND3_X1 \RegFile/_5859_ ( .A1(\RegFile/_1588_ ), .A2(\RegFile/_1527_ ), .A3(\RegFile/_3390_ ), .ZN(\RegFile/_1802_ ) );
NAND2_X1 \RegFile/_5860_ ( .A1(\RegFile/_1801_ ), .A2(\RegFile/_1802_ ), .ZN(\RegFile/_1803_ ) );
NOR4_X1 \RegFile/_5861_ ( .A1(\RegFile/_1798_ ), .A2(\RegFile/_1799_ ), .A3(\RegFile/_1800_ ), .A4(\RegFile/_1803_ ), .ZN(\RegFile/_1804_ ) );
NAND3_X1 \RegFile/_5862_ ( .A1(\RegFile/_1532_ ), .A2(\RegFile/_1536_ ), .A3(\RegFile/_3582_ ), .ZN(\RegFile/_1805_ ) );
INV_X1 \RegFile/_5863_ ( .A(\RegFile/_3614_ ), .ZN(\RegFile/_1806_ ) );
INV_X1 \RegFile/_5864_ ( .A(\RegFile/_3550_ ), .ZN(\RegFile/_1807_ ) );
OAI221_X1 \RegFile/_5865_ ( .A(\RegFile/_1805_ ), .B1(\RegFile/_1476_ ), .B2(\RegFile/_1806_ ), .C1(\RegFile/_1807_ ), .C2(\RegFile/_1512_ ), .ZN(\RegFile/_1808_ ) );
AND3_X1 \RegFile/_5866_ ( .A1(\RegFile/_1539_ ), .A2(\RegFile/_1429_ ), .A3(\RegFile/_3774_ ), .ZN(\RegFile/_1809_ ) );
NAND3_X1 \RegFile/_5867_ ( .A1(\RegFile/_1387_ ), .A2(\RegFile/_3742_ ), .A3(\RegFile/_1389_ ), .ZN(\RegFile/_1810_ ) );
OAI21_X1 \RegFile/_5868_ ( .A(\RegFile/_1810_ ), .B1(\RegFile/_1466_ ), .B2(\RegFile/_1187_ ), .ZN(\RegFile/_1811_ ) );
NOR4_X1 \RegFile/_5869_ ( .A1(\RegFile/_1808_ ), .A2(\RegFile/_1417_ ), .A3(\RegFile/_1809_ ), .A4(\RegFile/_1811_ ), .ZN(\RegFile/_1812_ ) );
BUF_X4 \RegFile/_5870_ ( .A(\RegFile/_1441_ ), .Z(\RegFile/_1813_ ) );
AOI22_X1 \RegFile/_5871_ ( .A1(\RegFile/_1804_ ), .A2(\RegFile/_1812_ ), .B1(\RegFile/_0086_ ), .B2(\RegFile/_1813_ ), .ZN(\RegFile/_0692_ ) );
NAND3_X1 \RegFile/_5872_ ( .A1(\RegFile/_1507_ ), .A2(\RegFile/_1472_ ), .A3(\RegFile/_3583_ ), .ZN(\RegFile/_1814_ ) );
INV_X1 \RegFile/_5873_ ( .A(\RegFile/_3615_ ), .ZN(\RegFile/_1815_ ) );
INV_X1 \RegFile/_5874_ ( .A(\RegFile/_3551_ ), .ZN(\RegFile/_1816_ ) );
OAI221_X1 \RegFile/_5875_ ( .A(\RegFile/_1814_ ), .B1(\RegFile/_1477_ ), .B2(\RegFile/_1815_ ), .C1(\RegFile/_1816_ ), .C2(\RegFile/_1512_ ), .ZN(\RegFile/_1817_ ) );
NAND3_X1 \RegFile/_5876_ ( .A1(\RegFile/_1468_ ), .A2(\RegFile/_3743_ ), .A3(\RegFile/_1484_ ), .ZN(\RegFile/_1818_ ) );
INV_X1 \RegFile/_5877_ ( .A(\RegFile/_3711_ ), .ZN(\RegFile/_1819_ ) );
OAI21_X1 \RegFile/_5878_ ( .A(\RegFile/_1818_ ), .B1(\RegFile/_1486_ ), .B2(\RegFile/_1819_ ), .ZN(\RegFile/_1820_ ) );
AND3_X1 \RegFile/_5879_ ( .A1(\RegFile/_1539_ ), .A2(\RegFile/_1558_ ), .A3(\RegFile/_3775_ ), .ZN(\RegFile/_1821_ ) );
NOR4_X1 \RegFile/_5880_ ( .A1(\RegFile/_1817_ ), .A2(\RegFile/_1480_ ), .A3(\RegFile/_1820_ ), .A4(\RegFile/_1821_ ), .ZN(\RegFile/_1822_ ) );
NAND3_X1 \RegFile/_5881_ ( .A1(\RegFile/_1420_ ), .A2(\RegFile/_1489_ ), .A3(\RegFile/_3679_ ), .ZN(\RegFile/_1823_ ) );
NAND3_X1 \RegFile/_5882_ ( .A1(\RegFile/_1393_ ), .A2(\RegFile/_3519_ ), .A3(\RegFile/_1396_ ), .ZN(\RegFile/_1824_ ) );
NAND3_X1 \RegFile/_5883_ ( .A1(\RegFile/_1443_ ), .A2(\RegFile/_1403_ ), .A3(\RegFile/_3327_ ), .ZN(\RegFile/_1825_ ) );
NAND3_X1 \RegFile/_5884_ ( .A1(\RegFile/_1443_ ), .A2(\RegFile/_3359_ ), .A3(\RegFile/_1421_ ), .ZN(\RegFile/_1826_ ) );
NAND3_X1 \RegFile/_5885_ ( .A1(\RegFile/_1431_ ), .A2(\RegFile/_1388_ ), .A3(\RegFile/_3391_ ), .ZN(\RegFile/_1827_ ) );
AND4_X1 \RegFile/_5886_ ( .A1(\RegFile/_1824_ ), .A2(\RegFile/_1825_ ), .A3(\RegFile/_1826_ ), .A4(\RegFile/_1827_ ), .ZN(\RegFile/_1828_ ) );
NAND3_X1 \RegFile/_5887_ ( .A1(\RegFile/_1430_ ), .A2(\RegFile/_3423_ ), .A3(\RegFile/_1526_ ), .ZN(\RegFile/_1829_ ) );
AOI22_X1 \RegFile/_5888_ ( .A1(\RegFile/_3647_ ), .A2(\RegFile/_1427_ ), .B1(\RegFile/_1407_ ), .B2(\RegFile/_1210_ ), .ZN(\RegFile/_1830_ ) );
AND4_X1 \RegFile/_5889_ ( .A1(\RegFile/_1823_ ), .A2(\RegFile/_1828_ ), .A3(\RegFile/_1829_ ), .A4(\RegFile/_1830_ ), .ZN(\RegFile/_1831_ ) );
AOI22_X1 \RegFile/_5890_ ( .A1(\RegFile/_1822_ ), .A2(\RegFile/_1831_ ), .B1(\RegFile/_0088_ ), .B2(\RegFile/_1813_ ), .ZN(\RegFile/_0693_ ) );
NAND3_X1 \RegFile/_5891_ ( .A1(\RegFile/_1471_ ), .A2(\RegFile/_3552_ ), .A3(\RegFile/_1508_ ), .ZN(\RegFile/_1832_ ) );
INV_X1 \RegFile/_5892_ ( .A(\RegFile/_3584_ ), .ZN(\RegFile/_1833_ ) );
INV_X1 \RegFile/_5893_ ( .A(\RegFile/_3616_ ), .ZN(\RegFile/_1834_ ) );
OAI221_X1 \RegFile/_5894_ ( .A(\RegFile/_1832_ ), .B1(\RegFile/_1474_ ), .B2(\RegFile/_1833_ ), .C1(\RegFile/_1477_ ), .C2(\RegFile/_1834_ ), .ZN(\RegFile/_1835_ ) );
AND3_X1 \RegFile/_5895_ ( .A1(\RegFile/_1481_ ), .A2(\RegFile/_1482_ ), .A3(\RegFile/_3776_ ), .ZN(\RegFile/_1836_ ) );
NAND3_X1 \RegFile/_5896_ ( .A1(\RegFile/_1468_ ), .A2(\RegFile/_3744_ ), .A3(\RegFile/_1464_ ), .ZN(\RegFile/_1837_ ) );
INV_X1 \RegFile/_5897_ ( .A(\RegFile/_3712_ ), .ZN(\RegFile/_1838_ ) );
OAI21_X1 \RegFile/_5898_ ( .A(\RegFile/_1837_ ), .B1(\RegFile/_1486_ ), .B2(\RegFile/_1838_ ), .ZN(\RegFile/_1839_ ) );
NOR4_X1 \RegFile/_5899_ ( .A1(\RegFile/_1835_ ), .A2(\RegFile/_1480_ ), .A3(\RegFile/_1836_ ), .A4(\RegFile/_1839_ ), .ZN(\RegFile/_1840_ ) );
NAND3_X1 \RegFile/_5900_ ( .A1(\RegFile/_1524_ ), .A2(\RegFile/_1577_ ), .A3(\RegFile/_3648_ ), .ZN(\RegFile/_1841_ ) );
NAND3_X1 \RegFile/_5901_ ( .A1(\RegFile/_1455_ ), .A2(\RegFile/_3424_ ), .A3(\RegFile/_1526_ ), .ZN(\RegFile/_1842_ ) );
NAND3_X1 \RegFile/_5902_ ( .A1(\RegFile/_1471_ ), .A2(\RegFile/_1226_ ), .A3(\RegFile/_1526_ ), .ZN(\RegFile/_1843_ ) );
NAND3_X1 \RegFile/_5903_ ( .A1(\RegFile/_1419_ ), .A2(\RegFile/_1530_ ), .A3(\RegFile/_3680_ ), .ZN(\RegFile/_1844_ ) );
NAND4_X1 \RegFile/_5904_ ( .A1(\RegFile/_1841_ ), .A2(\RegFile/_1842_ ), .A3(\RegFile/_1843_ ), .A4(\RegFile/_1844_ ), .ZN(\RegFile/_1845_ ) );
NAND3_X1 \RegFile/_5905_ ( .A1(\RegFile/_1583_ ), .A2(\RegFile/_1471_ ), .A3(\RegFile/_3328_ ), .ZN(\RegFile/_1846_ ) );
NAND3_X1 \RegFile/_5906_ ( .A1(\RegFile/_1529_ ), .A2(\RegFile/_3360_ ), .A3(\RegFile/_1532_ ), .ZN(\RegFile/_1847_ ) );
NAND2_X1 \RegFile/_5907_ ( .A1(\RegFile/_1846_ ), .A2(\RegFile/_1847_ ), .ZN(\RegFile/_1848_ ) );
AND3_X1 \RegFile/_5908_ ( .A1(\RegFile/_1482_ ), .A2(\RegFile/_3520_ ), .A3(\RegFile/_1536_ ), .ZN(\RegFile/_1849_ ) );
AND3_X1 \RegFile/_5909_ ( .A1(\RegFile/_1562_ ), .A2(\RegFile/_3392_ ), .A3(\RegFile/_1484_ ), .ZN(\RegFile/_1850_ ) );
NOR4_X1 \RegFile/_5910_ ( .A1(\RegFile/_1845_ ), .A2(\RegFile/_1848_ ), .A3(\RegFile/_1849_ ), .A4(\RegFile/_1850_ ), .ZN(\RegFile/_1851_ ) );
AOI22_X1 \RegFile/_5911_ ( .A1(\RegFile/_1840_ ), .A2(\RegFile/_1851_ ), .B1(\RegFile/_0090_ ), .B2(\RegFile/_1813_ ), .ZN(\RegFile/_0694_ ) );
NAND3_X1 \RegFile/_5912_ ( .A1(\RegFile/_1577_ ), .A2(\RegFile/_3617_ ), .A3(\RegFile/_1620_ ), .ZN(\RegFile/_1852_ ) );
INV_X1 \RegFile/_5913_ ( .A(\RegFile/_3585_ ), .ZN(\RegFile/_1853_ ) );
INV_X1 \RegFile/_5914_ ( .A(\RegFile/_3553_ ), .ZN(\RegFile/_1854_ ) );
OAI221_X1 \RegFile/_5915_ ( .A(\RegFile/_1852_ ), .B1(\RegFile/_1474_ ), .B2(\RegFile/_1853_ ), .C1(\RegFile/_1512_ ), .C2(\RegFile/_1854_ ), .ZN(\RegFile/_1855_ ) );
AND3_X1 \RegFile/_5916_ ( .A1(\RegFile/_1481_ ), .A2(\RegFile/_1482_ ), .A3(\RegFile/_3777_ ), .ZN(\RegFile/_1856_ ) );
NAND3_X1 \RegFile/_5917_ ( .A1(\RegFile/_1468_ ), .A2(\RegFile/_3745_ ), .A3(\RegFile/_1464_ ), .ZN(\RegFile/_1857_ ) );
INV_X1 \RegFile/_5918_ ( .A(\RegFile/_3713_ ), .ZN(\RegFile/_1858_ ) );
OAI21_X1 \RegFile/_5919_ ( .A(\RegFile/_1857_ ), .B1(\RegFile/_1466_ ), .B2(\RegFile/_1858_ ), .ZN(\RegFile/_1859_ ) );
NOR4_X1 \RegFile/_5920_ ( .A1(\RegFile/_1855_ ), .A2(\RegFile/_1441_ ), .A3(\RegFile/_1856_ ), .A4(\RegFile/_1859_ ), .ZN(\RegFile/_1860_ ) );
NAND3_X1 \RegFile/_5921_ ( .A1(\RegFile/_1420_ ), .A2(\RegFile/_1489_ ), .A3(\RegFile/_3681_ ), .ZN(\RegFile/_1861_ ) );
NAND3_X1 \RegFile/_5922_ ( .A1(\RegFile/_1393_ ), .A2(\RegFile/_3521_ ), .A3(\RegFile/_1396_ ), .ZN(\RegFile/_1862_ ) );
NAND3_X1 \RegFile/_5923_ ( .A1(\RegFile/_1443_ ), .A2(\RegFile/_1403_ ), .A3(\RegFile/_3329_ ), .ZN(\RegFile/_1863_ ) );
NAND3_X1 \RegFile/_5924_ ( .A1(\RegFile/_1443_ ), .A2(\RegFile/_3361_ ), .A3(\RegFile/_1421_ ), .ZN(\RegFile/_1864_ ) );
NAND3_X1 \RegFile/_5925_ ( .A1(\RegFile/_1431_ ), .A2(\RegFile/_1388_ ), .A3(\RegFile/_3393_ ), .ZN(\RegFile/_1865_ ) );
AND4_X1 \RegFile/_5926_ ( .A1(\RegFile/_1862_ ), .A2(\RegFile/_1863_ ), .A3(\RegFile/_1864_ ), .A4(\RegFile/_1865_ ), .ZN(\RegFile/_1866_ ) );
NAND3_X1 \RegFile/_5927_ ( .A1(\RegFile/_1430_ ), .A2(\RegFile/_3425_ ), .A3(\RegFile/_1526_ ), .ZN(\RegFile/_1867_ ) );
AOI22_X1 \RegFile/_5928_ ( .A1(\RegFile/_3649_ ), .A2(\RegFile/_1427_ ), .B1(\RegFile/_1407_ ), .B2(\RegFile/_1242_ ), .ZN(\RegFile/_1868_ ) );
AND4_X1 \RegFile/_5929_ ( .A1(\RegFile/_1861_ ), .A2(\RegFile/_1866_ ), .A3(\RegFile/_1867_ ), .A4(\RegFile/_1868_ ), .ZN(\RegFile/_1869_ ) );
AOI22_X1 \RegFile/_5930_ ( .A1(\RegFile/_1860_ ), .A2(\RegFile/_1869_ ), .B1(\RegFile/_0092_ ), .B2(\RegFile/_1813_ ), .ZN(\RegFile/_0695_ ) );
AND3_X1 \RegFile/_5931_ ( .A1(\RegFile/_1392_ ), .A2(\RegFile/_3522_ ), .A3(\RegFile/_1395_ ), .ZN(\RegFile/_1870_ ) );
NAND3_X1 \RegFile/_5932_ ( .A1(\RegFile/_1402_ ), .A2(\RegFile/_1258_ ), .A3(\RegFile/_1406_ ), .ZN(\RegFile/_1871_ ) );
OAI21_X1 \RegFile/_5933_ ( .A(\RegFile/_1871_ ), .B1(\RegFile/_1458_ ), .B2(\RegFile/_1248_ ), .ZN(\RegFile/_1872_ ) );
AOI211_X4 \RegFile/_5934_ ( .A(\RegFile/_1870_ ), .B(\RegFile/_1872_ ), .C1(\RegFile/_3554_ ), .C2(\RegFile/_1412_ ), .ZN(\RegFile/_1873_ ) );
AOI21_X1 \RegFile/_5935_ ( .A(\RegFile/_1416_ ), .B1(\RegFile/_1594_ ), .B2(\RegFile/_3778_ ), .ZN(\RegFile/_1874_ ) );
NAND3_X1 \RegFile/_5936_ ( .A1(\RegFile/_1596_ ), .A2(\RegFile/_3746_ ), .A3(\RegFile/_1434_ ), .ZN(\RegFile/_1875_ ) );
NAND3_X1 \RegFile/_5937_ ( .A1(\RegFile/_1430_ ), .A2(\RegFile/_1420_ ), .A3(\RegFile/_3650_ ), .ZN(\RegFile/_1876_ ) );
AND4_X1 \RegFile/_5938_ ( .A1(\RegFile/_1873_ ), .A2(\RegFile/_1874_ ), .A3(\RegFile/_1875_ ), .A4(\RegFile/_1876_ ), .ZN(\RegFile/_1877_ ) );
AND3_X1 \RegFile/_5939_ ( .A1(\RegFile/_1600_ ), .A2(\RegFile/_3586_ ), .A3(\RegFile/_1395_ ), .ZN(\RegFile/_1878_ ) );
AOI221_X4 \RegFile/_5940_ ( .A(\RegFile/_1878_ ), .B1(\RegFile/_1448_ ), .B2(\RegFile/_3618_ ), .C1(\RegFile/_3362_ ), .C2(\RegFile/_1437_ ), .ZN(\RegFile/_1879_ ) );
AOI22_X1 \RegFile/_5941_ ( .A1(\RegFile/_3330_ ), .A2(\RegFile/_1444_ ), .B1(\RegFile/_1461_ ), .B2(\RegFile/_3426_ ), .ZN(\RegFile/_1880_ ) );
NAND3_X1 \RegFile/_5942_ ( .A1(\RegFile/_1432_ ), .A2(\RegFile/_1620_ ), .A3(\RegFile/_3394_ ), .ZN(\RegFile/_1881_ ) );
NAND3_X1 \RegFile/_5943_ ( .A1(\RegFile/_1606_ ), .A2(\RegFile/_3714_ ), .A3(\RegFile/_1507_ ), .ZN(\RegFile/_1882_ ) );
AND4_X1 \RegFile/_5944_ ( .A1(\RegFile/_1879_ ), .A2(\RegFile/_1880_ ), .A3(\RegFile/_1881_ ), .A4(\RegFile/_1882_ ), .ZN(\RegFile/_1883_ ) );
AOI22_X1 \RegFile/_5945_ ( .A1(\RegFile/_1877_ ), .A2(\RegFile/_1883_ ), .B1(\RegFile/_0094_ ), .B2(\RegFile/_1813_ ), .ZN(\RegFile/_0696_ ) );
NOR2_X1 \RegFile/_5946_ ( .A1(\RegFile/_1409_ ), .A2(\RegFile/_0097_ ), .ZN(\RegFile/_1884_ ) );
AOI221_X4 \RegFile/_5947_ ( .A(\RegFile/_1884_ ), .B1(\RegFile/_3363_ ), .B2(\RegFile/_1437_ ), .C1(\RegFile/_3651_ ), .C2(\RegFile/_1427_ ), .ZN(\RegFile/_1885_ ) );
NAND3_X1 \RegFile/_5948_ ( .A1(\RegFile/_1596_ ), .A2(\RegFile/_1489_ ), .A3(\RegFile/_3331_ ), .ZN(\RegFile/_1886_ ) );
NAND3_X1 \RegFile/_5949_ ( .A1(\RegFile/_1489_ ), .A2(\RegFile/_3555_ ), .A3(\RegFile/_1472_ ), .ZN(\RegFile/_1887_ ) );
AOI22_X1 \RegFile/_5950_ ( .A1(\RegFile/_1426_ ), .A2(\RegFile/_3779_ ), .B1(\RegFile/_1451_ ), .B2(\RegFile/_3395_ ), .ZN(\RegFile/_1888_ ) );
AND4_X1 \RegFile/_5951_ ( .A1(\RegFile/_1885_ ), .A2(\RegFile/_1886_ ), .A3(\RegFile/_1887_ ), .A4(\RegFile/_1888_ ), .ZN(\RegFile/_1889_ ) );
AOI22_X1 \RegFile/_5952_ ( .A1(\RegFile/_1450_ ), .A2(\RegFile/_3523_ ), .B1(\RegFile/_1519_ ), .B2(\RegFile/_3683_ ), .ZN(\RegFile/_1890_ ) );
INV_X1 \RegFile/_5953_ ( .A(\RegFile/_3619_ ), .ZN(\RegFile/_1891_ ) );
OAI221_X1 \RegFile/_5954_ ( .A(\RegFile/_1890_ ), .B1(\RegFile/_1891_ ), .B2(\RegFile/_1476_ ), .C1(\RegFile/_1271_ ), .C2(\RegFile/_1474_ ), .ZN(\RegFile/_1892_ ) );
NAND4_X1 \RegFile/_5955_ ( .A1(\RegFile/_1389_ ), .A2(\RegFile/_3747_ ), .A3(\RegFile/_1384_ ), .A4(\RegFile/_0647_ ), .ZN(\RegFile/_1893_ ) );
OAI21_X1 \RegFile/_5956_ ( .A(\RegFile/_1893_ ), .B1(\RegFile/_1466_ ), .B2(\RegFile/_1275_ ), .ZN(\RegFile/_1894_ ) );
AND3_X1 \RegFile/_5957_ ( .A1(\RegFile/_1558_ ), .A2(\RegFile/_3427_ ), .A3(\RegFile/_1562_ ), .ZN(\RegFile/_1895_ ) );
NOR4_X1 \RegFile/_5958_ ( .A1(\RegFile/_1892_ ), .A2(\RegFile/_1417_ ), .A3(\RegFile/_1894_ ), .A4(\RegFile/_1895_ ), .ZN(\RegFile/_1896_ ) );
AOI22_X1 \RegFile/_5959_ ( .A1(\RegFile/_1889_ ), .A2(\RegFile/_1896_ ), .B1(\RegFile/_0096_ ), .B2(\RegFile/_1813_ ), .ZN(\RegFile/_0697_ ) );
AOI22_X1 \RegFile/_5960_ ( .A1(\RegFile/_3684_ ), .A2(\RegFile/_1519_ ), .B1(\RegFile/_1460_ ), .B2(\RegFile/_3428_ ), .ZN(\RegFile/_1897_ ) );
OAI221_X1 \RegFile/_5961_ ( .A(\RegFile/_1897_ ), .B1(\RegFile/_1521_ ), .B2(\RegFile/_0099_ ), .C1(\RegFile/_1281_ ), .C2(\RegFile/_1522_ ), .ZN(\RegFile/_1898_ ) );
AND3_X1 \RegFile/_5962_ ( .A1(\RegFile/_1455_ ), .A2(\RegFile/_3524_ ), .A3(\RegFile/_1508_ ), .ZN(\RegFile/_1899_ ) );
AND3_X1 \RegFile/_5963_ ( .A1(\RegFile/_1588_ ), .A2(\RegFile/_3396_ ), .A3(\RegFile/_1527_ ), .ZN(\RegFile/_1900_ ) );
NAND3_X1 \RegFile/_5964_ ( .A1(\RegFile/_1529_ ), .A2(\RegFile/_1530_ ), .A3(\RegFile/_3332_ ), .ZN(\RegFile/_1901_ ) );
NAND3_X1 \RegFile/_5965_ ( .A1(\RegFile/_1555_ ), .A2(\RegFile/_3364_ ), .A3(\RegFile/_1560_ ), .ZN(\RegFile/_1902_ ) );
NAND2_X1 \RegFile/_5966_ ( .A1(\RegFile/_1901_ ), .A2(\RegFile/_1902_ ), .ZN(\RegFile/_1903_ ) );
NOR4_X1 \RegFile/_5967_ ( .A1(\RegFile/_1898_ ), .A2(\RegFile/_1899_ ), .A3(\RegFile/_1900_ ), .A4(\RegFile/_1903_ ), .ZN(\RegFile/_1904_ ) );
AOI21_X1 \RegFile/_5968_ ( .A(\RegFile/_1417_ ), .B1(\RegFile/_1594_ ), .B2(\RegFile/_3780_ ), .ZN(\RegFile/_1905_ ) );
AND3_X1 \RegFile/_5969_ ( .A1(\RegFile/_1600_ ), .A2(\RegFile/_3588_ ), .A3(\RegFile/_1394_ ), .ZN(\RegFile/_1906_ ) );
AOI221_X4 \RegFile/_5970_ ( .A(\RegFile/_1906_ ), .B1(\RegFile/_1447_ ), .B2(\RegFile/_3620_ ), .C1(\RegFile/_3556_ ), .C2(\RegFile/_1411_ ), .ZN(\RegFile/_1907_ ) );
NAND3_X1 \RegFile/_5971_ ( .A1(\RegFile/_1583_ ), .A2(\RegFile/_3748_ ), .A3(\RegFile/_1620_ ), .ZN(\RegFile/_1908_ ) );
NAND3_X1 \RegFile/_5972_ ( .A1(\RegFile/_1606_ ), .A2(\RegFile/_3716_ ), .A3(\RegFile/_1507_ ), .ZN(\RegFile/_1909_ ) );
AND4_X1 \RegFile/_5973_ ( .A1(\RegFile/_1905_ ), .A2(\RegFile/_1907_ ), .A3(\RegFile/_1908_ ), .A4(\RegFile/_1909_ ), .ZN(\RegFile/_1910_ ) );
AOI22_X1 \RegFile/_5974_ ( .A1(\RegFile/_1904_ ), .A2(\RegFile/_1910_ ), .B1(\RegFile/_0098_ ), .B2(\RegFile/_1813_ ), .ZN(\RegFile/_0698_ ) );
NAND3_X1 \RegFile/_5975_ ( .A1(\RegFile/_1419_ ), .A2(\RegFile/_3621_ ), .A3(\RegFile/_1527_ ), .ZN(\RegFile/_1911_ ) );
INV_X1 \RegFile/_5976_ ( .A(\RegFile/_3589_ ), .ZN(\RegFile/_1912_ ) );
INV_X1 \RegFile/_5977_ ( .A(\RegFile/_3557_ ), .ZN(\RegFile/_1913_ ) );
OAI221_X1 \RegFile/_5978_ ( .A(\RegFile/_1911_ ), .B1(\RegFile/_1474_ ), .B2(\RegFile/_1912_ ), .C1(\RegFile/_1512_ ), .C2(\RegFile/_1913_ ), .ZN(\RegFile/_1914_ ) );
NAND3_X1 \RegFile/_5979_ ( .A1(\RegFile/_1468_ ), .A2(\RegFile/_3749_ ), .A3(\RegFile/_1484_ ), .ZN(\RegFile/_1915_ ) );
INV_X1 \RegFile/_5980_ ( .A(\RegFile/_3717_ ), .ZN(\RegFile/_1916_ ) );
OAI21_X1 \RegFile/_5981_ ( .A(\RegFile/_1915_ ), .B1(\RegFile/_1486_ ), .B2(\RegFile/_1916_ ), .ZN(\RegFile/_1917_ ) );
AND3_X1 \RegFile/_5982_ ( .A1(\RegFile/_1539_ ), .A2(\RegFile/_1558_ ), .A3(\RegFile/_3781_ ), .ZN(\RegFile/_1918_ ) );
NOR4_X1 \RegFile/_5983_ ( .A1(\RegFile/_1914_ ), .A2(\RegFile/_1441_ ), .A3(\RegFile/_1917_ ), .A4(\RegFile/_1918_ ), .ZN(\RegFile/_1919_ ) );
INV_X1 \RegFile/_5984_ ( .A(\RegFile/_3653_ ), .ZN(\RegFile/_1920_ ) );
OAI22_X1 \RegFile/_5985_ ( .A1(\RegFile/_1522_ ), .A2(\RegFile/_1920_ ), .B1(\RegFile/_1521_ ), .B2(\RegFile/_0101_ ), .ZN(\RegFile/_1921_ ) );
NAND3_X1 \RegFile/_5986_ ( .A1(\RegFile/_1555_ ), .A2(\RegFile/_1556_ ), .A3(\RegFile/_3333_ ), .ZN(\RegFile/_1922_ ) );
NAND3_X1 \RegFile/_5987_ ( .A1(\RegFile/_1429_ ), .A2(\RegFile/_3525_ ), .A3(\RegFile/_1396_ ), .ZN(\RegFile/_1923_ ) );
NAND3_X1 \RegFile/_5988_ ( .A1(\RegFile/_1387_ ), .A2(\RegFile/_3365_ ), .A3(\RegFile/_1560_ ), .ZN(\RegFile/_1924_ ) );
NAND3_X1 \RegFile/_5989_ ( .A1(\RegFile/_1562_ ), .A2(\RegFile/_1464_ ), .A3(\RegFile/_3397_ ), .ZN(\RegFile/_1925_ ) );
NAND4_X1 \RegFile/_5990_ ( .A1(\RegFile/_1922_ ), .A2(\RegFile/_1923_ ), .A3(\RegFile/_1924_ ), .A4(\RegFile/_1925_ ), .ZN(\RegFile/_1926_ ) );
AND3_X1 \RegFile/_5991_ ( .A1(\RegFile/_1419_ ), .A2(\RegFile/_1556_ ), .A3(\RegFile/_3685_ ), .ZN(\RegFile/_1927_ ) );
AND3_X1 \RegFile/_5992_ ( .A1(\RegFile/_1558_ ), .A2(\RegFile/_3429_ ), .A3(\RegFile/_1431_ ), .ZN(\RegFile/_1928_ ) );
NOR4_X1 \RegFile/_5993_ ( .A1(\RegFile/_1921_ ), .A2(\RegFile/_1926_ ), .A3(\RegFile/_1927_ ), .A4(\RegFile/_1928_ ), .ZN(\RegFile/_1929_ ) );
AOI22_X1 \RegFile/_5994_ ( .A1(\RegFile/_1919_ ), .A2(\RegFile/_1929_ ), .B1(\RegFile/_0100_ ), .B2(\RegFile/_1813_ ), .ZN(\RegFile/_0699_ ) );
AOI22_X1 \RegFile/_5995_ ( .A1(\RegFile/_3686_ ), .A2(\RegFile/_1519_ ), .B1(\RegFile/_1460_ ), .B2(\RegFile/_3430_ ), .ZN(\RegFile/_1930_ ) );
OAI221_X1 \RegFile/_5996_ ( .A(\RegFile/_1930_ ), .B1(\RegFile/_1521_ ), .B2(\RegFile/_0103_ ), .C1(\RegFile/_1315_ ), .C2(\RegFile/_1522_ ), .ZN(\RegFile/_1931_ ) );
AND3_X1 \RegFile/_5997_ ( .A1(\RegFile/_1455_ ), .A2(\RegFile/_3526_ ), .A3(\RegFile/_1508_ ), .ZN(\RegFile/_1932_ ) );
AND3_X1 \RegFile/_5998_ ( .A1(\RegFile/_1588_ ), .A2(\RegFile/_3398_ ), .A3(\RegFile/_1527_ ), .ZN(\RegFile/_1933_ ) );
NAND3_X1 \RegFile/_5999_ ( .A1(\RegFile/_1529_ ), .A2(\RegFile/_1530_ ), .A3(\RegFile/_3334_ ), .ZN(\RegFile/_1934_ ) );
NAND3_X1 \RegFile/_6000_ ( .A1(\RegFile/_1555_ ), .A2(\RegFile/_3366_ ), .A3(\RegFile/_1560_ ), .ZN(\RegFile/_1935_ ) );
NAND2_X1 \RegFile/_6001_ ( .A1(\RegFile/_1934_ ), .A2(\RegFile/_1935_ ), .ZN(\RegFile/_1936_ ) );
NOR4_X1 \RegFile/_6002_ ( .A1(\RegFile/_1931_ ), .A2(\RegFile/_1932_ ), .A3(\RegFile/_1933_ ), .A4(\RegFile/_1936_ ), .ZN(\RegFile/_1937_ ) );
AOI21_X1 \RegFile/_6003_ ( .A(\RegFile/_1417_ ), .B1(\RegFile/_1594_ ), .B2(\RegFile/_3782_ ), .ZN(\RegFile/_1938_ ) );
AND3_X1 \RegFile/_6004_ ( .A1(\RegFile/_1414_ ), .A2(\RegFile/_3590_ ), .A3(\RegFile/_1394_ ), .ZN(\RegFile/_1939_ ) );
AOI221_X4 \RegFile/_6005_ ( .A(\RegFile/_1939_ ), .B1(\RegFile/_1447_ ), .B2(\RegFile/_3622_ ), .C1(\RegFile/_3558_ ), .C2(\RegFile/_1411_ ), .ZN(\RegFile/_1940_ ) );
NAND3_X1 \RegFile/_6006_ ( .A1(\RegFile/_1583_ ), .A2(\RegFile/_3750_ ), .A3(\RegFile/_1620_ ), .ZN(\RegFile/_1941_ ) );
NAND3_X1 \RegFile/_6007_ ( .A1(\RegFile/_1606_ ), .A2(\RegFile/_3718_ ), .A3(\RegFile/_1507_ ), .ZN(\RegFile/_1942_ ) );
AND4_X1 \RegFile/_6008_ ( .A1(\RegFile/_1938_ ), .A2(\RegFile/_1940_ ), .A3(\RegFile/_1941_ ), .A4(\RegFile/_1942_ ), .ZN(\RegFile/_1943_ ) );
AOI22_X1 \RegFile/_6009_ ( .A1(\RegFile/_1937_ ), .A2(\RegFile/_1943_ ), .B1(\RegFile/_0102_ ), .B2(\RegFile/_1813_ ), .ZN(\RegFile/_0700_ ) );
NAND3_X1 \RegFile/_6010_ ( .A1(\RegFile/_1596_ ), .A2(\RegFile/_3751_ ), .A3(\RegFile/_1434_ ), .ZN(\RegFile/_1944_ ) );
AND3_X1 \RegFile/_6011_ ( .A1(\RegFile/_1600_ ), .A2(\RegFile/_3591_ ), .A3(\RegFile/_1394_ ), .ZN(\RegFile/_1945_ ) );
AOI221_X4 \RegFile/_6012_ ( .A(\RegFile/_1945_ ), .B1(\RegFile/_1448_ ), .B2(\RegFile/_3623_ ), .C1(\RegFile/_3559_ ), .C2(\RegFile/_1412_ ), .ZN(\RegFile/_1946_ ) );
NAND3_X1 \RegFile/_6013_ ( .A1(\RegFile/_1420_ ), .A2(\RegFile/_3719_ ), .A3(\RegFile/_1422_ ), .ZN(\RegFile/_1947_ ) );
AOI21_X1 \RegFile/_6014_ ( .A(\RegFile/_1416_ ), .B1(\RegFile/_1426_ ), .B2(\RegFile/_3783_ ), .ZN(\RegFile/_1948_ ) );
AND4_X1 \RegFile/_6015_ ( .A1(\RegFile/_1944_ ), .A2(\RegFile/_1946_ ), .A3(\RegFile/_1947_ ), .A4(\RegFile/_1948_ ), .ZN(\RegFile/_1949_ ) );
NAND3_X1 \RegFile/_6016_ ( .A1(\RegFile/_1489_ ), .A2(\RegFile/_1345_ ), .A3(\RegFile/_1432_ ), .ZN(\RegFile/_1950_ ) );
AOI22_X1 \RegFile/_6017_ ( .A1(\RegFile/_3687_ ), .A2(\RegFile/_1519_ ), .B1(\RegFile/_1461_ ), .B2(\RegFile/_3431_ ), .ZN(\RegFile/_1951_ ) );
NAND3_X1 \RegFile/_6018_ ( .A1(\RegFile/_1393_ ), .A2(\RegFile/_3527_ ), .A3(\RegFile/_1396_ ), .ZN(\RegFile/_1952_ ) );
NAND3_X1 \RegFile/_6019_ ( .A1(\RegFile/_1443_ ), .A2(\RegFile/_1403_ ), .A3(\RegFile/_3335_ ), .ZN(\RegFile/_1953_ ) );
NAND3_X1 \RegFile/_6020_ ( .A1(\RegFile/_1386_ ), .A2(\RegFile/_3367_ ), .A3(\RegFile/_1421_ ), .ZN(\RegFile/_1954_ ) );
NAND3_X1 \RegFile/_6021_ ( .A1(\RegFile/_1431_ ), .A2(\RegFile/_1388_ ), .A3(\RegFile/_3399_ ), .ZN(\RegFile/_1955_ ) );
AND4_X1 \RegFile/_6022_ ( .A1(\RegFile/_1952_ ), .A2(\RegFile/_1953_ ), .A3(\RegFile/_1954_ ), .A4(\RegFile/_1955_ ), .ZN(\RegFile/_1956_ ) );
NAND3_X1 \RegFile/_6023_ ( .A1(\RegFile/_1524_ ), .A2(\RegFile/_1577_ ), .A3(\RegFile/_3655_ ), .ZN(\RegFile/_1957_ ) );
AND4_X1 \RegFile/_6024_ ( .A1(\RegFile/_1950_ ), .A2(\RegFile/_1951_ ), .A3(\RegFile/_1956_ ), .A4(\RegFile/_1957_ ), .ZN(\RegFile/_1958_ ) );
AOI22_X1 \RegFile/_6025_ ( .A1(\RegFile/_1949_ ), .A2(\RegFile/_1958_ ), .B1(\RegFile/_0104_ ), .B2(\RegFile/_1813_ ), .ZN(\RegFile/_0701_ ) );
AOI22_X1 \RegFile/_6026_ ( .A1(\RegFile/_3689_ ), .A2(\RegFile/_1519_ ), .B1(\RegFile/_1460_ ), .B2(\RegFile/_3433_ ), .ZN(\RegFile/_1959_ ) );
OAI221_X1 \RegFile/_6027_ ( .A(\RegFile/_1959_ ), .B1(\RegFile/_1409_ ), .B2(\RegFile/_0107_ ), .C1(\RegFile/_1353_ ), .C2(\RegFile/_1500_ ), .ZN(\RegFile/_1960_ ) );
AND3_X1 \RegFile/_6028_ ( .A1(\RegFile/_1455_ ), .A2(\RegFile/_3529_ ), .A3(\RegFile/_1508_ ), .ZN(\RegFile/_1961_ ) );
AND3_X1 \RegFile/_6029_ ( .A1(\RegFile/_1588_ ), .A2(\RegFile/_3401_ ), .A3(\RegFile/_1527_ ), .ZN(\RegFile/_1962_ ) );
NAND3_X1 \RegFile/_6030_ ( .A1(\RegFile/_1481_ ), .A2(\RegFile/_1556_ ), .A3(\RegFile/_3337_ ), .ZN(\RegFile/_1963_ ) );
NAND3_X1 \RegFile/_6031_ ( .A1(\RegFile/_1555_ ), .A2(\RegFile/_3369_ ), .A3(\RegFile/_1560_ ), .ZN(\RegFile/_1964_ ) );
NAND2_X1 \RegFile/_6032_ ( .A1(\RegFile/_1963_ ), .A2(\RegFile/_1964_ ), .ZN(\RegFile/_1965_ ) );
NOR4_X1 \RegFile/_6033_ ( .A1(\RegFile/_1960_ ), .A2(\RegFile/_1961_ ), .A3(\RegFile/_1962_ ), .A4(\RegFile/_1965_ ), .ZN(\RegFile/_1966_ ) );
AOI21_X1 \RegFile/_6034_ ( .A(\RegFile/_1416_ ), .B1(\RegFile/_1594_ ), .B2(\RegFile/_3785_ ), .ZN(\RegFile/_1967_ ) );
AND3_X1 \RegFile/_6035_ ( .A1(\RegFile/_1414_ ), .A2(\RegFile/_3593_ ), .A3(\RegFile/_1394_ ), .ZN(\RegFile/_1968_ ) );
AOI221_X4 \RegFile/_6036_ ( .A(\RegFile/_1968_ ), .B1(\RegFile/_1447_ ), .B2(\RegFile/_3625_ ), .C1(\RegFile/_3561_ ), .C2(\RegFile/_1411_ ), .ZN(\RegFile/_1969_ ) );
NAND3_X1 \RegFile/_6037_ ( .A1(\RegFile/_1583_ ), .A2(\RegFile/_3753_ ), .A3(\RegFile/_1620_ ), .ZN(\RegFile/_1970_ ) );
NAND3_X1 \RegFile/_6038_ ( .A1(\RegFile/_1606_ ), .A2(\RegFile/_3721_ ), .A3(\RegFile/_1507_ ), .ZN(\RegFile/_1971_ ) );
AND4_X1 \RegFile/_6039_ ( .A1(\RegFile/_1967_ ), .A2(\RegFile/_1969_ ), .A3(\RegFile/_1970_ ), .A4(\RegFile/_1971_ ), .ZN(\RegFile/_1972_ ) );
AOI22_X1 \RegFile/_6040_ ( .A1(\RegFile/_1966_ ), .A2(\RegFile/_1972_ ), .B1(\RegFile/_0106_ ), .B2(\RegFile/_1480_ ), .ZN(\RegFile/_0703_ ) );
NAND3_X1 \RegFile/_6041_ ( .A1(\RegFile/_1399_ ), .A2(\RegFile/_1402_ ), .A3(\RegFile/_3690_ ), .ZN(\RegFile/_1973_ ) );
OAI21_X1 \RegFile/_6042_ ( .A(\RegFile/_1973_ ), .B1(\RegFile/_1409_ ), .B2(\RegFile/_0109_ ), .ZN(\RegFile/_1974_ ) );
AOI221_X4 \RegFile/_6043_ ( .A(\RegFile/_1974_ ), .B1(\RegFile/_3562_ ), .B2(\RegFile/_1411_ ), .C1(\RegFile/_3530_ ), .C2(\RegFile/_1450_ ), .ZN(\RegFile/_1975_ ) );
AOI21_X1 \RegFile/_6044_ ( .A(\RegFile/_1416_ ), .B1(\RegFile/_1594_ ), .B2(\RegFile/_3786_ ), .ZN(\RegFile/_1976_ ) );
NAND3_X1 \RegFile/_6045_ ( .A1(\RegFile/_1596_ ), .A2(\RegFile/_3754_ ), .A3(\RegFile/_1434_ ), .ZN(\RegFile/_1977_ ) );
NAND3_X1 \RegFile/_6046_ ( .A1(\RegFile/_1430_ ), .A2(\RegFile/_1606_ ), .A3(\RegFile/_3658_ ), .ZN(\RegFile/_1978_ ) );
AND4_X1 \RegFile/_6047_ ( .A1(\RegFile/_1975_ ), .A2(\RegFile/_1976_ ), .A3(\RegFile/_1977_ ), .A4(\RegFile/_1978_ ), .ZN(\RegFile/_1979_ ) );
AND3_X1 \RegFile/_6048_ ( .A1(\RegFile/_1600_ ), .A2(\RegFile/_3594_ ), .A3(\RegFile/_1395_ ), .ZN(\RegFile/_1980_ ) );
AOI221_X4 \RegFile/_6049_ ( .A(\RegFile/_1980_ ), .B1(\RegFile/_1448_ ), .B2(\RegFile/_3626_ ), .C1(\RegFile/_3370_ ), .C2(\RegFile/_1437_ ), .ZN(\RegFile/_1981_ ) );
AND3_X1 \RegFile/_6050_ ( .A1(\RegFile/_1386_ ), .A2(\RegFile/_1402_ ), .A3(\RegFile/_3338_ ), .ZN(\RegFile/_1982_ ) );
AOI21_X1 \RegFile/_6051_ ( .A(\RegFile/_1982_ ), .B1(\RegFile/_3434_ ), .B2(\RegFile/_1461_ ), .ZN(\RegFile/_1983_ ) );
NAND3_X1 \RegFile/_6052_ ( .A1(\RegFile/_1432_ ), .A2(\RegFile/_1620_ ), .A3(\RegFile/_3402_ ), .ZN(\RegFile/_1984_ ) );
NAND3_X1 \RegFile/_6053_ ( .A1(\RegFile/_1577_ ), .A2(\RegFile/_3722_ ), .A3(\RegFile/_1507_ ), .ZN(\RegFile/_1985_ ) );
AND4_X1 \RegFile/_6054_ ( .A1(\RegFile/_1981_ ), .A2(\RegFile/_1983_ ), .A3(\RegFile/_1984_ ), .A4(\RegFile/_1985_ ), .ZN(\RegFile/_1986_ ) );
AOI22_X1 \RegFile/_6055_ ( .A1(\RegFile/_1979_ ), .A2(\RegFile/_1986_ ), .B1(\RegFile/_0108_ ), .B2(\RegFile/_1480_ ), .ZN(\RegFile/_0704_ ) );
AND2_X4 \RegFile/_6056_ ( .A1(\RegFile/_0713_ ), .A2(\RegFile/_0712_ ), .ZN(\RegFile/_1987_ ) );
BUF_X8 \RegFile/_6057_ ( .A(\RegFile/_1987_ ), .Z(\RegFile/_1988_ ) );
BUF_X4 \RegFile/_6058_ ( .A(\RegFile/_1988_ ), .Z(\RegFile/_1989_ ) );
BUF_X4 \RegFile/_6059_ ( .A(\RegFile/_1989_ ), .Z(\RegFile/_1990_ ) );
BUF_X4 \RegFile/_6060_ ( .A(\RegFile/_1990_ ), .Z(\RegFile/_1991_ ) );
AND2_X4 \RegFile/_6061_ ( .A1(\RegFile/_0715_ ), .A2(\RegFile/_0714_ ), .ZN(\RegFile/_1992_ ) );
BUF_X8 \RegFile/_6062_ ( .A(\RegFile/_1992_ ), .Z(\RegFile/_1993_ ) );
BUF_X16 \RegFile/_6063_ ( .A(\RegFile/_1993_ ), .Z(\RegFile/_1994_ ) );
BUF_X4 \RegFile/_6064_ ( .A(\RegFile/_1994_ ), .Z(\RegFile/_1995_ ) );
BUF_X4 \RegFile/_6065_ ( .A(\RegFile/_1995_ ), .Z(\RegFile/_1996_ ) );
BUF_X4 \RegFile/_6066_ ( .A(\RegFile/_1996_ ), .Z(\RegFile/_1997_ ) );
AOI21_X1 \RegFile/_6067_ ( .A(\RegFile/_3474_ ), .B1(\RegFile/_1991_ ), .B2(\RegFile/_1997_ ), .ZN(\RegFile/_1998_ ) );
INV_X16 \RegFile/_6068_ ( .A(\RegFile/_0714_ ), .ZN(\RegFile/_1999_ ) );
AND2_X4 \RegFile/_6069_ ( .A1(\RegFile/_1999_ ), .A2(\RegFile/_0715_ ), .ZN(\RegFile/_2000_ ) );
BUF_X8 \RegFile/_6070_ ( .A(\RegFile/_2000_ ), .Z(\RegFile/_2001_ ) );
NOR2_X4 \RegFile/_6071_ ( .A1(\RegFile/_0713_ ), .A2(\RegFile/_0712_ ), .ZN(\RegFile/_2002_ ) );
BUF_X4 \RegFile/_6072_ ( .A(\RegFile/_2002_ ), .Z(\RegFile/_2003_ ) );
AND2_X2 \RegFile/_6073_ ( .A1(\RegFile/_2001_ ), .A2(\RegFile/_2003_ ), .ZN(\RegFile/_2004_ ) );
BUF_X4 \RegFile/_6074_ ( .A(\RegFile/_2004_ ), .Z(\RegFile/_2005_ ) );
NOR2_X4 \RegFile/_6075_ ( .A1(\RegFile/_1999_ ), .A2(\RegFile/_0715_ ), .ZN(\RegFile/_2006_ ) );
AND2_X1 \RegFile/_6076_ ( .A1(\RegFile/_2006_ ), .A2(\RegFile/_1987_ ), .ZN(\RegFile/_2007_ ) );
BUF_X4 \RegFile/_6077_ ( .A(\RegFile/_2007_ ), .Z(\RegFile/_2008_ ) );
BUF_X4 \RegFile/_6078_ ( .A(\RegFile/_2008_ ), .Z(\RegFile/_2009_ ) );
AOI22_X1 \RegFile/_6079_ ( .A1(\RegFile/_2005_ ), .A2(\RegFile/_3730_ ), .B1(\RegFile/_2009_ ), .B2(\RegFile/_3698_ ), .ZN(\RegFile/_2010_ ) );
INV_X32 \RegFile/_6080_ ( .A(\RegFile/_0713_ ), .ZN(\RegFile/_2011_ ) );
AND2_X4 \RegFile/_6081_ ( .A1(\RegFile/_2011_ ), .A2(\RegFile/_0712_ ), .ZN(\RegFile/_2012_ ) );
AND2_X1 \RegFile/_6082_ ( .A1(\RegFile/_2001_ ), .A2(\RegFile/_2012_ ), .ZN(\RegFile/_2013_ ) );
BUF_X4 \RegFile/_6083_ ( .A(\RegFile/_2013_ ), .Z(\RegFile/_2014_ ) );
NOR2_X1 \RegFile/_6084_ ( .A1(\RegFile/_2011_ ), .A2(\RegFile/_0712_ ), .ZN(\RegFile/_2015_ ) );
AND2_X1 \RegFile/_6085_ ( .A1(\RegFile/_2000_ ), .A2(\RegFile/_2015_ ), .ZN(\RegFile/_2016_ ) );
BUF_X4 \RegFile/_6086_ ( .A(\RegFile/_2016_ ), .Z(\RegFile/_2017_ ) );
BUF_X4 \RegFile/_6087_ ( .A(\RegFile/_2017_ ), .Z(\RegFile/_2018_ ) );
AOI22_X1 \RegFile/_6088_ ( .A1(\RegFile/_3762_ ), .A2(\RegFile/_2014_ ), .B1(\RegFile/_2018_ ), .B2(\RegFile/_3314_ ), .ZN(\RegFile/_2019_ ) );
AND2_X2 \RegFile/_6089_ ( .A1(\RegFile/_2001_ ), .A2(\RegFile/_1987_ ), .ZN(\RegFile/_2020_ ) );
BUF_X4 \RegFile/_6090_ ( .A(\RegFile/_2020_ ), .Z(\RegFile/_2021_ ) );
AND2_X4 \RegFile/_6091_ ( .A1(\RegFile/_1993_ ), .A2(\RegFile/_2002_ ), .ZN(\RegFile/_2022_ ) );
BUF_X4 \RegFile/_6092_ ( .A(\RegFile/_2022_ ), .Z(\RegFile/_2023_ ) );
BUF_X4 \RegFile/_6093_ ( .A(\RegFile/_2023_ ), .Z(\RegFile/_2024_ ) );
AOI22_X1 \RegFile/_6094_ ( .A1(\RegFile/_2021_ ), .A2(\RegFile/_3346_ ), .B1(\RegFile/_3378_ ), .B2(\RegFile/_2024_ ), .ZN(\RegFile/_2025_ ) );
BUF_X4 \RegFile/_6095_ ( .A(\RegFile/_2015_ ), .Z(\RegFile/_2026_ ) );
BUF_X2 \RegFile/_6096_ ( .A(\RegFile/_2026_ ), .Z(\RegFile/_2027_ ) );
BUF_X4 \RegFile/_6097_ ( .A(\RegFile/_1993_ ), .Z(\RegFile/_2028_ ) );
AND3_X1 \RegFile/_6098_ ( .A1(\RegFile/_2027_ ), .A2(\RegFile/_3442_ ), .A3(\RegFile/_2028_ ), .ZN(\RegFile/_2029_ ) );
AND2_X2 \RegFile/_6099_ ( .A1(\RegFile/_2012_ ), .A2(\RegFile/_1993_ ), .ZN(\RegFile/_2030_ ) );
BUF_X4 \RegFile/_6100_ ( .A(\RegFile/_2030_ ), .Z(\RegFile/_2031_ ) );
AOI21_X1 \RegFile/_6101_ ( .A(\RegFile/_2029_ ), .B1(\RegFile/_3410_ ), .B2(\RegFile/_2031_ ), .ZN(\RegFile/_2032_ ) );
AND4_X1 \RegFile/_6102_ ( .A1(\RegFile/_2010_ ), .A2(\RegFile/_2019_ ), .A3(\RegFile/_2025_ ), .A4(\RegFile/_2032_ ), .ZN(\RegFile/_2033_ ) );
BUF_X4 \RegFile/_6103_ ( .A(\RegFile/_2003_ ), .Z(\RegFile/_2034_ ) );
BUF_X4 \RegFile/_6104_ ( .A(\RegFile/_2034_ ), .Z(\RegFile/_2035_ ) );
NOR2_X4 \RegFile/_6105_ ( .A1(\RegFile/_0715_ ), .A2(\RegFile/_0714_ ), .ZN(\RegFile/_2036_ ) );
BUF_X4 \RegFile/_6106_ ( .A(\RegFile/_2036_ ), .Z(\RegFile/_2037_ ) );
BUF_X4 \RegFile/_6107_ ( .A(\RegFile/_2037_ ), .Z(\RegFile/_2038_ ) );
NAND3_X1 \RegFile/_6108_ ( .A1(\RegFile/_2035_ ), .A2(\RegFile/_2038_ ), .A3(\RegFile/_3282_ ), .ZN(\RegFile/_2039_ ) );
CLKBUF_X2 \RegFile/_6109_ ( .A(\RegFile/_2006_ ), .Z(\RegFile/_2040_ ) );
BUF_X2 \RegFile/_6110_ ( .A(\RegFile/_2026_ ), .Z(\RegFile/_2041_ ) );
AND3_X1 \RegFile/_6111_ ( .A1(\RegFile/_2040_ ), .A2(\RegFile/_2041_ ), .A3(\RegFile/_3666_ ), .ZN(\RegFile/_2042_ ) );
AND2_X2 \RegFile/_6112_ ( .A1(\RegFile/_2012_ ), .A2(\RegFile/_2006_ ), .ZN(\RegFile/_2043_ ) );
BUF_X4 \RegFile/_6113_ ( .A(\RegFile/_2043_ ), .Z(\RegFile/_2044_ ) );
BUF_X4 \RegFile/_6114_ ( .A(\RegFile/_2044_ ), .Z(\RegFile/_2045_ ) );
AOI21_X1 \RegFile/_6115_ ( .A(\RegFile/_2042_ ), .B1(\RegFile/_3634_ ), .B2(\RegFile/_2045_ ), .ZN(\RegFile/_2046_ ) );
AND2_X2 \RegFile/_6116_ ( .A1(\RegFile/_2012_ ), .A2(\RegFile/_2037_ ), .ZN(\RegFile/_2047_ ) );
BUF_X4 \RegFile/_6117_ ( .A(\RegFile/_2047_ ), .Z(\RegFile/_2048_ ) );
AND2_X2 \RegFile/_6118_ ( .A1(\RegFile/_2015_ ), .A2(\RegFile/_2037_ ), .ZN(\RegFile/_2049_ ) );
BUF_X4 \RegFile/_6119_ ( .A(\RegFile/_2049_ ), .Z(\RegFile/_2050_ ) );
AOI22_X1 \RegFile/_6120_ ( .A1(\RegFile/_2048_ ), .A2(\RegFile/_3506_ ), .B1(\RegFile/_2050_ ), .B2(\RegFile/_3538_ ), .ZN(\RegFile/_2051_ ) );
AND2_X2 \RegFile/_6121_ ( .A1(\RegFile/_2006_ ), .A2(\RegFile/_2003_ ), .ZN(\RegFile/_2052_ ) );
BUF_X4 \RegFile/_6122_ ( .A(\RegFile/_2052_ ), .Z(\RegFile/_2053_ ) );
AND2_X2 \RegFile/_6123_ ( .A1(\RegFile/_1987_ ), .A2(\RegFile/_2036_ ), .ZN(\RegFile/_2054_ ) );
BUF_X4 \RegFile/_6124_ ( .A(\RegFile/_2054_ ), .Z(\RegFile/_2055_ ) );
AOI22_X1 \RegFile/_6125_ ( .A1(\RegFile/_2053_ ), .A2(\RegFile/_3602_ ), .B1(\RegFile/_2055_ ), .B2(\RegFile/_3570_ ), .ZN(\RegFile/_2056_ ) );
AND4_X1 \RegFile/_6126_ ( .A1(\RegFile/_2039_ ), .A2(\RegFile/_2046_ ), .A3(\RegFile/_2051_ ), .A4(\RegFile/_2056_ ), .ZN(\RegFile/_2057_ ) );
AND2_X4 \RegFile/_6127_ ( .A1(\RegFile/_2002_ ), .A2(\RegFile/_2037_ ), .ZN(\RegFile/_2058_ ) );
BUF_X8 \RegFile/_6128_ ( .A(\RegFile/_2058_ ), .Z(\RegFile/_2059_ ) );
INV_X1 \RegFile/_6129_ ( .A(\RegFile/_0748_ ), .ZN(\RegFile/_2060_ ) );
NOR2_X2 \RegFile/_6130_ ( .A1(\RegFile/_2059_ ), .A2(\RegFile/_2060_ ), .ZN(\RegFile/_2061_ ) );
INV_X2 \RegFile/_6131_ ( .A(\RegFile/_2061_ ), .ZN(\RegFile/_2062_ ) );
BUF_X4 \RegFile/_6132_ ( .A(\RegFile/_2062_ ), .Z(\RegFile/_2063_ ) );
NAND3_X1 \RegFile/_6133_ ( .A1(\RegFile/_1990_ ), .A2(\RegFile/_1996_ ), .A3(\RegFile/_3474_ ), .ZN(\RegFile/_2064_ ) );
NAND4_X1 \RegFile/_6134_ ( .A1(\RegFile/_2033_ ), .A2(\RegFile/_2057_ ), .A3(\RegFile/_2063_ ), .A4(\RegFile/_2064_ ), .ZN(\RegFile/_2065_ ) );
BUF_X2 \RegFile/_6135_ ( .A(\RegFile/_2059_ ), .Z(\RegFile/_2066_ ) );
BUF_X2 \RegFile/_6136_ ( .A(\RegFile/_2066_ ), .Z(\RegFile/_2067_ ) );
BUF_X2 \RegFile/_6137_ ( .A(\RegFile/_2060_ ), .Z(\RegFile/_2068_ ) );
BUF_X2 \RegFile/_6138_ ( .A(\RegFile/_2068_ ), .Z(\RegFile/_2069_ ) );
OR3_X1 \RegFile/_6139_ ( .A1(\RegFile/_2067_ ), .A2(\RegFile/_2069_ ), .A3(\RegFile/_0716_ ), .ZN(\RegFile/_2070_ ) );
NAND2_X1 \RegFile/_6140_ ( .A1(\RegFile/_2065_ ), .A2(\RegFile/_2070_ ), .ZN(\RegFile/_2071_ ) );
BUF_X4 \RegFile/_6141_ ( .A(\RegFile/_2071_ ), .Z(\RegFile/_2072_ ) );
AND2_X1 \RegFile/_6142_ ( .A1(\RegFile/_1987_ ), .A2(\RegFile/_1993_ ), .ZN(\RegFile/_2073_ ) );
BUF_X4 \RegFile/_6143_ ( .A(\RegFile/_2073_ ), .Z(\RegFile/_2074_ ) );
BUF_X4 \RegFile/_6144_ ( .A(\RegFile/_2074_ ), .Z(\RegFile/_2075_ ) );
AOI21_X1 \RegFile/_6145_ ( .A(\RegFile/_1998_ ), .B1(\RegFile/_2072_ ), .B2(\RegFile/_2075_ ), .ZN(\RegFile/_0608_ ) );
INV_X1 \RegFile/_6146_ ( .A(\RegFile/_2074_ ), .ZN(\RegFile/_2076_ ) );
BUF_X4 \RegFile/_6147_ ( .A(\RegFile/_2076_ ), .Z(\RegFile/_2077_ ) );
NAND2_X1 \RegFile/_6148_ ( .A1(\RegFile/_2077_ ), .A2(\RegFile/_3485_ ), .ZN(\RegFile/_2078_ ) );
AND3_X1 \RegFile/_6149_ ( .A1(\RegFile/_2040_ ), .A2(\RegFile/_2027_ ), .A3(\RegFile/_3677_ ), .ZN(\RegFile/_2079_ ) );
AOI21_X1 \RegFile/_6150_ ( .A(\RegFile/_2079_ ), .B1(\RegFile/_3709_ ), .B2(\RegFile/_2009_ ), .ZN(\RegFile/_2080_ ) );
BUF_X4 \RegFile/_6151_ ( .A(\RegFile/_2020_ ), .Z(\RegFile/_2081_ ) );
AOI22_X1 \RegFile/_6152_ ( .A1(\RegFile/_3325_ ), .A2(\RegFile/_2018_ ), .B1(\RegFile/_2081_ ), .B2(\RegFile/_3357_ ), .ZN(\RegFile/_2082_ ) );
BUF_X16 \RegFile/_6153_ ( .A(\RegFile/_2059_ ), .Z(\RegFile/_2083_ ) );
AOI22_X1 \RegFile/_6154_ ( .A1(\RegFile/_2048_ ), .A2(\RegFile/_3517_ ), .B1(\RegFile/_3293_ ), .B2(\RegFile/_2083_ ), .ZN(\RegFile/_2084_ ) );
BUF_X4 \RegFile/_6155_ ( .A(\RegFile/_2030_ ), .Z(\RegFile/_2085_ ) );
BUF_X4 \RegFile/_6156_ ( .A(\RegFile/_2022_ ), .Z(\RegFile/_2086_ ) );
AOI22_X1 \RegFile/_6157_ ( .A1(\RegFile/_2085_ ), .A2(\RegFile/_3421_ ), .B1(\RegFile/_3389_ ), .B2(\RegFile/_2086_ ), .ZN(\RegFile/_2087_ ) );
AND4_X1 \RegFile/_6158_ ( .A1(\RegFile/_2080_ ), .A2(\RegFile/_2082_ ), .A3(\RegFile/_2084_ ), .A4(\RegFile/_2087_ ), .ZN(\RegFile/_2088_ ) );
BUF_X4 \RegFile/_6159_ ( .A(\RegFile/_2062_ ), .Z(\RegFile/_2089_ ) );
CLKBUF_X2 \RegFile/_6160_ ( .A(\RegFile/_2015_ ), .Z(\RegFile/_2090_ ) );
BUF_X4 \RegFile/_6161_ ( .A(\RegFile/_2037_ ), .Z(\RegFile/_2091_ ) );
NAND3_X1 \RegFile/_6162_ ( .A1(\RegFile/_2090_ ), .A2(\RegFile/_3549_ ), .A3(\RegFile/_2091_ ), .ZN(\RegFile/_2092_ ) );
NAND3_X1 \RegFile/_6163_ ( .A1(\RegFile/_1988_ ), .A2(\RegFile/_2037_ ), .A3(\RegFile/_3581_ ), .ZN(\RegFile/_2093_ ) );
NAND2_X1 \RegFile/_6164_ ( .A1(\RegFile/_2092_ ), .A2(\RegFile/_2093_ ), .ZN(\RegFile/_2094_ ) );
AOI221_X4 \RegFile/_6165_ ( .A(\RegFile/_2094_ ), .B1(\RegFile/_3645_ ), .B2(\RegFile/_2044_ ), .C1(\RegFile/_3613_ ), .C2(\RegFile/_2053_ ), .ZN(\RegFile/_2095_ ) );
BUF_X4 \RegFile/_6166_ ( .A(\RegFile/_2001_ ), .Z(\RegFile/_2096_ ) );
BUF_X4 \RegFile/_6167_ ( .A(\RegFile/_2012_ ), .Z(\RegFile/_2097_ ) );
BUF_X4 \RegFile/_6168_ ( .A(\RegFile/_2097_ ), .Z(\RegFile/_2098_ ) );
NAND3_X1 \RegFile/_6169_ ( .A1(\RegFile/_2096_ ), .A2(\RegFile/_2098_ ), .A3(\RegFile/_3773_ ), .ZN(\RegFile/_2099_ ) );
BUF_X4 \RegFile/_6170_ ( .A(\RegFile/_2001_ ), .Z(\RegFile/_2100_ ) );
BUF_X4 \RegFile/_6171_ ( .A(\RegFile/_2003_ ), .Z(\RegFile/_2101_ ) );
NAND3_X1 \RegFile/_6172_ ( .A1(\RegFile/_2100_ ), .A2(\RegFile/_3741_ ), .A3(\RegFile/_2101_ ), .ZN(\RegFile/_2102_ ) );
BUF_X4 \RegFile/_6173_ ( .A(\RegFile/_1993_ ), .Z(\RegFile/_2103_ ) );
BUF_X4 \RegFile/_6174_ ( .A(\RegFile/_2103_ ), .Z(\RegFile/_2104_ ) );
NAND3_X1 \RegFile/_6175_ ( .A1(\RegFile/_1989_ ), .A2(\RegFile/_2104_ ), .A3(\RegFile/_3485_ ), .ZN(\RegFile/_2105_ ) );
BUF_X2 \RegFile/_6176_ ( .A(\RegFile/_2015_ ), .Z(\RegFile/_2106_ ) );
BUF_X4 \RegFile/_6177_ ( .A(\RegFile/_2106_ ), .Z(\RegFile/_2107_ ) );
NAND3_X1 \RegFile/_6178_ ( .A1(\RegFile/_2107_ ), .A2(\RegFile/_3453_ ), .A3(\RegFile/_2104_ ), .ZN(\RegFile/_2108_ ) );
AND4_X1 \RegFile/_6179_ ( .A1(\RegFile/_2099_ ), .A2(\RegFile/_2102_ ), .A3(\RegFile/_2105_ ), .A4(\RegFile/_2108_ ), .ZN(\RegFile/_2109_ ) );
NAND4_X1 \RegFile/_6180_ ( .A1(\RegFile/_2088_ ), .A2(\RegFile/_2089_ ), .A3(\RegFile/_2095_ ), .A4(\RegFile/_2109_ ), .ZN(\RegFile/_2110_ ) );
OR3_X1 \RegFile/_6181_ ( .A1(\RegFile/_2066_ ), .A2(\RegFile/_2068_ ), .A3(\RegFile/_0727_ ), .ZN(\RegFile/_2111_ ) );
NAND2_X1 \RegFile/_6182_ ( .A1(\RegFile/_2110_ ), .A2(\RegFile/_2111_ ), .ZN(\RegFile/_2112_ ) );
BUF_X4 \RegFile/_6183_ ( .A(\RegFile/_2112_ ), .Z(\RegFile/_2113_ ) );
BUF_X4 \RegFile/_6184_ ( .A(\RegFile/_2076_ ), .Z(\RegFile/_2114_ ) );
OAI21_X1 \RegFile/_6185_ ( .A(\RegFile/_2078_ ), .B1(\RegFile/_2113_ ), .B2(\RegFile/_2114_ ), .ZN(\RegFile/_0609_ ) );
NAND2_X1 \RegFile/_6186_ ( .A1(\RegFile/_2077_ ), .A2(\RegFile/_3496_ ), .ZN(\RegFile/_2115_ ) );
INV_X1 \RegFile/_6187_ ( .A(\RegFile/_2007_ ), .ZN(\RegFile/_2116_ ) );
BUF_X2 \RegFile/_6188_ ( .A(\RegFile/_2006_ ), .Z(\RegFile/_2117_ ) );
NAND2_X2 \RegFile/_6189_ ( .A1(\RegFile/_2117_ ), .A2(\RegFile/_2026_ ), .ZN(\RegFile/_2118_ ) );
OAI22_X1 \RegFile/_6190_ ( .A1(\RegFile/_2116_ ), .A2(\RegFile/_0859_ ), .B1(\RegFile/_2118_ ), .B2(\RegFile/_0856_ ), .ZN(\RegFile/_2119_ ) );
BUF_X4 \RegFile/_6191_ ( .A(\RegFile/_2047_ ), .Z(\RegFile/_2120_ ) );
BUF_X4 \RegFile/_6192_ ( .A(\RegFile/_2059_ ), .Z(\RegFile/_2121_ ) );
AOI221_X4 \RegFile/_6193_ ( .A(\RegFile/_2119_ ), .B1(\RegFile/_3528_ ), .B2(\RegFile/_2120_ ), .C1(\RegFile/_3304_ ), .C2(\RegFile/_2121_ ), .ZN(\RegFile/_2122_ ) );
NAND3_X1 \RegFile/_6194_ ( .A1(\RegFile/_2097_ ), .A2(\RegFile/_3432_ ), .A3(\RegFile/_1994_ ), .ZN(\RegFile/_2123_ ) );
NAND3_X1 \RegFile/_6195_ ( .A1(\RegFile/_2103_ ), .A2(\RegFile/_2003_ ), .A3(\RegFile/_3400_ ), .ZN(\RegFile/_2124_ ) );
NAND2_X1 \RegFile/_6196_ ( .A1(\RegFile/_2123_ ), .A2(\RegFile/_2124_ ), .ZN(\RegFile/_2125_ ) );
BUF_X4 \RegFile/_6197_ ( .A(\RegFile/_2020_ ), .Z(\RegFile/_2126_ ) );
BUF_X4 \RegFile/_6198_ ( .A(\RegFile/_2017_ ), .Z(\RegFile/_2127_ ) );
AOI221_X4 \RegFile/_6199_ ( .A(\RegFile/_2125_ ), .B1(\RegFile/_3368_ ), .B2(\RegFile/_2126_ ), .C1(\RegFile/_3336_ ), .C2(\RegFile/_2127_ ), .ZN(\RegFile/_2128_ ) );
AOI22_X1 \RegFile/_6200_ ( .A1(\RegFile/_2050_ ), .A2(\RegFile/_3560_ ), .B1(\RegFile/_2055_ ), .B2(\RegFile/_3592_ ), .ZN(\RegFile/_2129_ ) );
BUF_X4 \RegFile/_6201_ ( .A(\RegFile/_2013_ ), .Z(\RegFile/_2130_ ) );
BUF_X4 \RegFile/_6202_ ( .A(\RegFile/_2004_ ), .Z(\RegFile/_2131_ ) );
AOI22_X1 \RegFile/_6203_ ( .A1(\RegFile/_3784_ ), .A2(\RegFile/_2130_ ), .B1(\RegFile/_2131_ ), .B2(\RegFile/_3752_ ), .ZN(\RegFile/_2132_ ) );
BUF_X4 \RegFile/_6204_ ( .A(\RegFile/_2044_ ), .Z(\RegFile/_2133_ ) );
BUF_X4 \RegFile/_6205_ ( .A(\RegFile/_2052_ ), .Z(\RegFile/_2134_ ) );
AOI22_X1 \RegFile/_6206_ ( .A1(\RegFile/_2133_ ), .A2(\RegFile/_3656_ ), .B1(\RegFile/_2134_ ), .B2(\RegFile/_3624_ ), .ZN(\RegFile/_2135_ ) );
AND3_X1 \RegFile/_6207_ ( .A1(\RegFile/_2090_ ), .A2(\RegFile/_3464_ ), .A3(\RegFile/_1994_ ), .ZN(\RegFile/_2136_ ) );
AOI21_X1 \RegFile/_6208_ ( .A(\RegFile/_2136_ ), .B1(\RegFile/_3496_ ), .B2(\RegFile/_2074_ ), .ZN(\RegFile/_2137_ ) );
AND4_X1 \RegFile/_6209_ ( .A1(\RegFile/_2129_ ), .A2(\RegFile/_2132_ ), .A3(\RegFile/_2135_ ), .A4(\RegFile/_2137_ ), .ZN(\RegFile/_2138_ ) );
NAND4_X4 \RegFile/_6210_ ( .A1(\RegFile/_2122_ ), .A2(\RegFile/_2089_ ), .A3(\RegFile/_2128_ ), .A4(\RegFile/_2138_ ), .ZN(\RegFile/_2139_ ) );
OR3_X1 \RegFile/_6211_ ( .A1(\RegFile/_2066_ ), .A2(\RegFile/_2068_ ), .A3(\RegFile/_0738_ ), .ZN(\RegFile/_2140_ ) );
NAND2_X1 \RegFile/_6212_ ( .A1(\RegFile/_2139_ ), .A2(\RegFile/_2140_ ), .ZN(\RegFile/_2141_ ) );
BUF_X4 \RegFile/_6213_ ( .A(\RegFile/_2141_ ), .Z(\RegFile/_2142_ ) );
OAI21_X1 \RegFile/_6214_ ( .A(\RegFile/_2115_ ), .B1(\RegFile/_2142_ ), .B2(\RegFile/_2114_ ), .ZN(\RegFile/_0610_ ) );
AOI21_X1 \RegFile/_6215_ ( .A(\RegFile/_3499_ ), .B1(\RegFile/_1991_ ), .B2(\RegFile/_1997_ ), .ZN(\RegFile/_2143_ ) );
INV_X4 \RegFile/_6216_ ( .A(\RegFile/_2049_ ), .ZN(\RegFile/_2144_ ) );
INV_X4 \RegFile/_6217_ ( .A(\RegFile/_2054_ ), .ZN(\RegFile/_2145_ ) );
BUF_X4 \RegFile/_6218_ ( .A(\RegFile/_2145_ ), .Z(\RegFile/_2146_ ) );
INV_X1 \RegFile/_6219_ ( .A(\RegFile/_3595_ ), .ZN(\RegFile/_2147_ ) );
OAI22_X1 \RegFile/_6220_ ( .A1(\RegFile/_2144_ ), .A2(\RegFile/_1511_ ), .B1(\RegFile/_2146_ ), .B2(\RegFile/_2147_ ), .ZN(\RegFile/_2148_ ) );
BUF_X4 \RegFile/_6221_ ( .A(\RegFile/_2134_ ), .Z(\RegFile/_2149_ ) );
AOI221_X4 \RegFile/_6222_ ( .A(\RegFile/_2148_ ), .B1(\RegFile/_3659_ ), .B2(\RegFile/_2133_ ), .C1(\RegFile/_3627_ ), .C2(\RegFile/_2149_ ), .ZN(\RegFile/_2150_ ) );
AND3_X1 \RegFile/_6223_ ( .A1(\RegFile/_2040_ ), .A2(\RegFile/_2027_ ), .A3(\RegFile/_3691_ ), .ZN(\RegFile/_2151_ ) );
BUF_X4 \RegFile/_6224_ ( .A(\RegFile/_2008_ ), .Z(\RegFile/_2152_ ) );
AOI21_X1 \RegFile/_6225_ ( .A(\RegFile/_2151_ ), .B1(\RegFile/_3723_ ), .B2(\RegFile/_2152_ ), .ZN(\RegFile/_2153_ ) );
AOI22_X1 \RegFile/_6226_ ( .A1(\RegFile/_3339_ ), .A2(\RegFile/_2018_ ), .B1(\RegFile/_2081_ ), .B2(\RegFile/_3371_ ), .ZN(\RegFile/_2154_ ) );
BUF_X4 \RegFile/_6227_ ( .A(\RegFile/_2047_ ), .Z(\RegFile/_2155_ ) );
AOI22_X1 \RegFile/_6228_ ( .A1(\RegFile/_2155_ ), .A2(\RegFile/_3531_ ), .B1(\RegFile/_3307_ ), .B2(\RegFile/_2121_ ), .ZN(\RegFile/_2156_ ) );
AOI22_X1 \RegFile/_6229_ ( .A1(\RegFile/_2031_ ), .A2(\RegFile/_3435_ ), .B1(\RegFile/_3403_ ), .B2(\RegFile/_2024_ ), .ZN(\RegFile/_2157_ ) );
AND4_X1 \RegFile/_6230_ ( .A1(\RegFile/_2153_ ), .A2(\RegFile/_2154_ ), .A3(\RegFile/_2156_ ), .A4(\RegFile/_2157_ ), .ZN(\RegFile/_2158_ ) );
BUF_X4 \RegFile/_6231_ ( .A(\RegFile/_2001_ ), .Z(\RegFile/_2159_ ) );
BUF_X4 \RegFile/_6232_ ( .A(\RegFile/_2159_ ), .Z(\RegFile/_2160_ ) );
BUF_X4 \RegFile/_6233_ ( .A(\RegFile/_2097_ ), .Z(\RegFile/_2161_ ) );
NAND3_X1 \RegFile/_6234_ ( .A1(\RegFile/_2160_ ), .A2(\RegFile/_2161_ ), .A3(\RegFile/_3787_ ), .ZN(\RegFile/_2162_ ) );
BUF_X4 \RegFile/_6235_ ( .A(\RegFile/_2034_ ), .Z(\RegFile/_2163_ ) );
NAND3_X1 \RegFile/_6236_ ( .A1(\RegFile/_2096_ ), .A2(\RegFile/_3755_ ), .A3(\RegFile/_2163_ ), .ZN(\RegFile/_2164_ ) );
BUF_X4 \RegFile/_6237_ ( .A(\RegFile/_1988_ ), .Z(\RegFile/_2165_ ) );
BUF_X4 \RegFile/_6238_ ( .A(\RegFile/_2165_ ), .Z(\RegFile/_2166_ ) );
NAND3_X1 \RegFile/_6239_ ( .A1(\RegFile/_2166_ ), .A2(\RegFile/_1996_ ), .A3(\RegFile/_3499_ ), .ZN(\RegFile/_2167_ ) );
BUF_X4 \RegFile/_6240_ ( .A(\RegFile/_2026_ ), .Z(\RegFile/_2168_ ) );
BUF_X4 \RegFile/_6241_ ( .A(\RegFile/_2168_ ), .Z(\RegFile/_2169_ ) );
BUF_X4 \RegFile/_6242_ ( .A(\RegFile/_2028_ ), .Z(\RegFile/_2170_ ) );
NAND3_X1 \RegFile/_6243_ ( .A1(\RegFile/_2169_ ), .A2(\RegFile/_3467_ ), .A3(\RegFile/_2170_ ), .ZN(\RegFile/_2171_ ) );
AND4_X1 \RegFile/_6244_ ( .A1(\RegFile/_2162_ ), .A2(\RegFile/_2164_ ), .A3(\RegFile/_2167_ ), .A4(\RegFile/_2171_ ), .ZN(\RegFile/_2172_ ) );
NAND4_X4 \RegFile/_6245_ ( .A1(\RegFile/_2150_ ), .A2(\RegFile/_2063_ ), .A3(\RegFile/_2158_ ), .A4(\RegFile/_2172_ ), .ZN(\RegFile/_2173_ ) );
OR3_X2 \RegFile/_6246_ ( .A1(\RegFile/_2067_ ), .A2(\RegFile/_2069_ ), .A3(\RegFile/_0741_ ), .ZN(\RegFile/_2174_ ) );
NAND2_X2 \RegFile/_6247_ ( .A1(\RegFile/_2173_ ), .A2(\RegFile/_2174_ ), .ZN(\RegFile/_2175_ ) );
AOI21_X1 \RegFile/_6248_ ( .A(\RegFile/_2143_ ), .B1(\RegFile/_2175_ ), .B2(\RegFile/_2075_ ), .ZN(\RegFile/_0611_ ) );
AOI21_X1 \RegFile/_6249_ ( .A(\RegFile/_3500_ ), .B1(\RegFile/_1991_ ), .B2(\RegFile/_1997_ ), .ZN(\RegFile/_2176_ ) );
BUF_X4 \RegFile/_6250_ ( .A(\RegFile/_2054_ ), .Z(\RegFile/_2177_ ) );
AOI22_X1 \RegFile/_6251_ ( .A1(\RegFile/_2050_ ), .A2(\RegFile/_3564_ ), .B1(\RegFile/_2177_ ), .B2(\RegFile/_3596_ ), .ZN(\RegFile/_2178_ ) );
INV_X2 \RegFile/_6252_ ( .A(\RegFile/_2052_ ), .ZN(\RegFile/_2179_ ) );
BUF_X4 \RegFile/_6253_ ( .A(\RegFile/_2179_ ), .Z(\RegFile/_2180_ ) );
INV_X4 \RegFile/_6254_ ( .A(\RegFile/_2044_ ), .ZN(\RegFile/_2181_ ) );
BUF_X4 \RegFile/_6255_ ( .A(\RegFile/_2181_ ), .Z(\RegFile/_2182_ ) );
OAI221_X1 \RegFile/_6256_ ( .A(\RegFile/_2178_ ), .B1(\RegFile/_0910_ ), .B2(\RegFile/_2180_ ), .C1(\RegFile/_0902_ ), .C2(\RegFile/_2182_ ), .ZN(\RegFile/_2183_ ) );
AOI22_X1 \RegFile/_6257_ ( .A1(\RegFile/_3340_ ), .A2(\RegFile/_2017_ ), .B1(\RegFile/_2126_ ), .B2(\RegFile/_3372_ ), .ZN(\RegFile/_2184_ ) );
AND3_X1 \RegFile/_6258_ ( .A1(\RegFile/_2117_ ), .A2(\RegFile/_2026_ ), .A3(\RegFile/_3692_ ), .ZN(\RegFile/_2185_ ) );
AOI21_X1 \RegFile/_6259_ ( .A(\RegFile/_2185_ ), .B1(\RegFile/_3724_ ), .B2(\RegFile/_2008_ ), .ZN(\RegFile/_2186_ ) );
AOI22_X1 \RegFile/_6260_ ( .A1(\RegFile/_2120_ ), .A2(\RegFile/_3532_ ), .B1(\RegFile/_3308_ ), .B2(\RegFile/_2059_ ), .ZN(\RegFile/_2187_ ) );
BUF_X4 \RegFile/_6261_ ( .A(\RegFile/_2030_ ), .Z(\RegFile/_2188_ ) );
AOI22_X1 \RegFile/_6262_ ( .A1(\RegFile/_2188_ ), .A2(\RegFile/_3436_ ), .B1(\RegFile/_3404_ ), .B2(\RegFile/_2023_ ), .ZN(\RegFile/_2189_ ) );
NAND4_X1 \RegFile/_6263_ ( .A1(\RegFile/_2184_ ), .A2(\RegFile/_2186_ ), .A3(\RegFile/_2187_ ), .A4(\RegFile/_2189_ ), .ZN(\RegFile/_2190_ ) );
NAND3_X1 \RegFile/_6264_ ( .A1(\RegFile/_2100_ ), .A2(\RegFile/_2098_ ), .A3(\RegFile/_3788_ ), .ZN(\RegFile/_2191_ ) );
NAND3_X1 \RegFile/_6265_ ( .A1(\RegFile/_2100_ ), .A2(\RegFile/_3756_ ), .A3(\RegFile/_2101_ ), .ZN(\RegFile/_2192_ ) );
NAND3_X1 \RegFile/_6266_ ( .A1(\RegFile/_2165_ ), .A2(\RegFile/_1995_ ), .A3(\RegFile/_3500_ ), .ZN(\RegFile/_2193_ ) );
NAND3_X1 \RegFile/_6267_ ( .A1(\RegFile/_2107_ ), .A2(\RegFile/_3468_ ), .A3(\RegFile/_1995_ ), .ZN(\RegFile/_2194_ ) );
NAND4_X1 \RegFile/_6268_ ( .A1(\RegFile/_2191_ ), .A2(\RegFile/_2192_ ), .A3(\RegFile/_2193_ ), .A4(\RegFile/_2194_ ), .ZN(\RegFile/_2195_ ) );
NOR4_X1 \RegFile/_6269_ ( .A1(\RegFile/_2183_ ), .A2(\RegFile/_2190_ ), .A3(\RegFile/_2061_ ), .A4(\RegFile/_2195_ ), .ZN(\RegFile/_2196_ ) );
AOI211_X4 \RegFile/_6270_ ( .A(\RegFile/_2068_ ), .B(\RegFile/_0742_ ), .C1(\RegFile/_2035_ ), .C2(\RegFile/_2038_ ), .ZN(\RegFile/_2197_ ) );
OR2_X2 \RegFile/_6271_ ( .A1(\RegFile/_2196_ ), .A2(\RegFile/_2197_ ), .ZN(\RegFile/_2198_ ) );
BUF_X4 \RegFile/_6272_ ( .A(\RegFile/_2198_ ), .Z(\RegFile/_2199_ ) );
AOI21_X1 \RegFile/_6273_ ( .A(\RegFile/_2176_ ), .B1(\RegFile/_2199_ ), .B2(\RegFile/_2075_ ), .ZN(\RegFile/_0612_ ) );
AOI21_X1 \RegFile/_6274_ ( .A(\RegFile/_3501_ ), .B1(\RegFile/_1991_ ), .B2(\RegFile/_1997_ ), .ZN(\RegFile/_2200_ ) );
INV_X1 \RegFile/_6275_ ( .A(\RegFile/_3597_ ), .ZN(\RegFile/_2201_ ) );
OAI22_X1 \RegFile/_6276_ ( .A1(\RegFile/_2144_ ), .A2(\RegFile/_1546_ ), .B1(\RegFile/_2146_ ), .B2(\RegFile/_2201_ ), .ZN(\RegFile/_2202_ ) );
AOI221_X4 \RegFile/_6277_ ( .A(\RegFile/_2202_ ), .B1(\RegFile/_3661_ ), .B2(\RegFile/_2045_ ), .C1(\RegFile/_3629_ ), .C2(\RegFile/_2149_ ), .ZN(\RegFile/_2203_ ) );
AND3_X1 \RegFile/_6278_ ( .A1(\RegFile/_2040_ ), .A2(\RegFile/_2168_ ), .A3(\RegFile/_3693_ ), .ZN(\RegFile/_2204_ ) );
AOI21_X1 \RegFile/_6279_ ( .A(\RegFile/_2204_ ), .B1(\RegFile/_3725_ ), .B2(\RegFile/_2152_ ), .ZN(\RegFile/_2205_ ) );
BUF_X4 \RegFile/_6280_ ( .A(\RegFile/_2017_ ), .Z(\RegFile/_2206_ ) );
AOI22_X1 \RegFile/_6281_ ( .A1(\RegFile/_3341_ ), .A2(\RegFile/_2206_ ), .B1(\RegFile/_2021_ ), .B2(\RegFile/_3373_ ), .ZN(\RegFile/_2207_ ) );
AOI22_X1 \RegFile/_6282_ ( .A1(\RegFile/_2155_ ), .A2(\RegFile/_3533_ ), .B1(\RegFile/_3309_ ), .B2(\RegFile/_2121_ ), .ZN(\RegFile/_2208_ ) );
AOI22_X1 \RegFile/_6283_ ( .A1(\RegFile/_2031_ ), .A2(\RegFile/_3437_ ), .B1(\RegFile/_3405_ ), .B2(\RegFile/_2024_ ), .ZN(\RegFile/_2209_ ) );
AND4_X1 \RegFile/_6284_ ( .A1(\RegFile/_2205_ ), .A2(\RegFile/_2207_ ), .A3(\RegFile/_2208_ ), .A4(\RegFile/_2209_ ), .ZN(\RegFile/_2210_ ) );
NAND3_X1 \RegFile/_6285_ ( .A1(\RegFile/_2160_ ), .A2(\RegFile/_2161_ ), .A3(\RegFile/_3789_ ), .ZN(\RegFile/_2211_ ) );
NAND3_X1 \RegFile/_6286_ ( .A1(\RegFile/_2160_ ), .A2(\RegFile/_3757_ ), .A3(\RegFile/_2163_ ), .ZN(\RegFile/_2212_ ) );
NAND3_X1 \RegFile/_6287_ ( .A1(\RegFile/_2166_ ), .A2(\RegFile/_1996_ ), .A3(\RegFile/_3501_ ), .ZN(\RegFile/_2213_ ) );
NAND3_X1 \RegFile/_6288_ ( .A1(\RegFile/_2169_ ), .A2(\RegFile/_3469_ ), .A3(\RegFile/_2170_ ), .ZN(\RegFile/_2214_ ) );
AND4_X1 \RegFile/_6289_ ( .A1(\RegFile/_2211_ ), .A2(\RegFile/_2212_ ), .A3(\RegFile/_2213_ ), .A4(\RegFile/_2214_ ), .ZN(\RegFile/_2215_ ) );
NAND4_X4 \RegFile/_6290_ ( .A1(\RegFile/_2203_ ), .A2(\RegFile/_2063_ ), .A3(\RegFile/_2210_ ), .A4(\RegFile/_2215_ ), .ZN(\RegFile/_2216_ ) );
OR3_X2 \RegFile/_6291_ ( .A1(\RegFile/_2067_ ), .A2(\RegFile/_2069_ ), .A3(\RegFile/_0743_ ), .ZN(\RegFile/_2217_ ) );
NAND2_X2 \RegFile/_6292_ ( .A1(\RegFile/_2216_ ), .A2(\RegFile/_2217_ ), .ZN(\RegFile/_2218_ ) );
AOI21_X1 \RegFile/_6293_ ( .A(\RegFile/_2200_ ), .B1(\RegFile/_2218_ ), .B2(\RegFile/_2075_ ), .ZN(\RegFile/_0613_ ) );
AOI21_X1 \RegFile/_6294_ ( .A(\RegFile/_3502_ ), .B1(\RegFile/_1991_ ), .B2(\RegFile/_1997_ ), .ZN(\RegFile/_2219_ ) );
CLKBUF_X2 \RegFile/_6295_ ( .A(\RegFile/_2006_ ), .Z(\RegFile/_2220_ ) );
NAND3_X1 \RegFile/_6296_ ( .A1(\RegFile/_2220_ ), .A2(\RegFile/_2106_ ), .A3(\RegFile/_3694_ ), .ZN(\RegFile/_2221_ ) );
OAI21_X1 \RegFile/_6297_ ( .A(\RegFile/_2221_ ), .B1(\RegFile/_2116_ ), .B2(\RegFile/_1574_ ), .ZN(\RegFile/_2222_ ) );
AOI221_X4 \RegFile/_6298_ ( .A(\RegFile/_2222_ ), .B1(\RegFile/_3534_ ), .B2(\RegFile/_2120_ ), .C1(\RegFile/_3310_ ), .C2(\RegFile/_2066_ ), .ZN(\RegFile/_2223_ ) );
NAND3_X1 \RegFile/_6299_ ( .A1(\RegFile/_2097_ ), .A2(\RegFile/_3438_ ), .A3(\RegFile/_2103_ ), .ZN(\RegFile/_2224_ ) );
NAND3_X1 \RegFile/_6300_ ( .A1(\RegFile/_2103_ ), .A2(\RegFile/_2003_ ), .A3(\RegFile/_3406_ ), .ZN(\RegFile/_2225_ ) );
NAND2_X1 \RegFile/_6301_ ( .A1(\RegFile/_2224_ ), .A2(\RegFile/_2225_ ), .ZN(\RegFile/_2226_ ) );
AOI221_X4 \RegFile/_6302_ ( .A(\RegFile/_2226_ ), .B1(\RegFile/_3374_ ), .B2(\RegFile/_2126_ ), .C1(\RegFile/_3342_ ), .C2(\RegFile/_2127_ ), .ZN(\RegFile/_2227_ ) );
BUF_X4 \RegFile/_6303_ ( .A(\RegFile/_2049_ ), .Z(\RegFile/_2228_ ) );
AOI22_X1 \RegFile/_6304_ ( .A1(\RegFile/_2228_ ), .A2(\RegFile/_3566_ ), .B1(\RegFile/_2055_ ), .B2(\RegFile/_3598_ ), .ZN(\RegFile/_2229_ ) );
AOI22_X1 \RegFile/_6305_ ( .A1(\RegFile/_3790_ ), .A2(\RegFile/_2130_ ), .B1(\RegFile/_2131_ ), .B2(\RegFile/_3758_ ), .ZN(\RegFile/_2230_ ) );
AOI22_X1 \RegFile/_6306_ ( .A1(\RegFile/_2133_ ), .A2(\RegFile/_3662_ ), .B1(\RegFile/_2134_ ), .B2(\RegFile/_3630_ ), .ZN(\RegFile/_2231_ ) );
AND3_X1 \RegFile/_6307_ ( .A1(\RegFile/_2090_ ), .A2(\RegFile/_3470_ ), .A3(\RegFile/_1994_ ), .ZN(\RegFile/_2232_ ) );
AOI21_X1 \RegFile/_6308_ ( .A(\RegFile/_2232_ ), .B1(\RegFile/_3502_ ), .B2(\RegFile/_2074_ ), .ZN(\RegFile/_2233_ ) );
AND4_X1 \RegFile/_6309_ ( .A1(\RegFile/_2229_ ), .A2(\RegFile/_2230_ ), .A3(\RegFile/_2231_ ), .A4(\RegFile/_2233_ ), .ZN(\RegFile/_2234_ ) );
NAND4_X4 \RegFile/_6310_ ( .A1(\RegFile/_2223_ ), .A2(\RegFile/_2089_ ), .A3(\RegFile/_2227_ ), .A4(\RegFile/_2234_ ), .ZN(\RegFile/_2235_ ) );
CLKBUF_X2 \RegFile/_6311_ ( .A(\RegFile/_2066_ ), .Z(\RegFile/_2236_ ) );
CLKBUF_X2 \RegFile/_6312_ ( .A(\RegFile/_2068_ ), .Z(\RegFile/_2237_ ) );
OR3_X1 \RegFile/_6313_ ( .A1(\RegFile/_2236_ ), .A2(\RegFile/_2237_ ), .A3(\RegFile/_0744_ ), .ZN(\RegFile/_2238_ ) );
NAND2_X1 \RegFile/_6314_ ( .A1(\RegFile/_2235_ ), .A2(\RegFile/_2238_ ), .ZN(\RegFile/_2239_ ) );
BUF_X4 \RegFile/_6315_ ( .A(\RegFile/_2239_ ), .Z(\RegFile/_2240_ ) );
AOI21_X1 \RegFile/_6316_ ( .A(\RegFile/_2219_ ), .B1(\RegFile/_2240_ ), .B2(\RegFile/_2075_ ), .ZN(\RegFile/_0614_ ) );
AOI21_X1 \RegFile/_6317_ ( .A(\RegFile/_3503_ ), .B1(\RegFile/_1991_ ), .B2(\RegFile/_1997_ ), .ZN(\RegFile/_2241_ ) );
NAND3_X1 \RegFile/_6318_ ( .A1(\RegFile/_2220_ ), .A2(\RegFile/_3631_ ), .A3(\RegFile/_2034_ ), .ZN(\RegFile/_2242_ ) );
OAI21_X1 \RegFile/_6319_ ( .A(\RegFile/_2242_ ), .B1(\RegFile/_2182_ ), .B2(\RegFile/_0959_ ), .ZN(\RegFile/_2243_ ) );
AOI221_X1 \RegFile/_6320_ ( .A(\RegFile/_2243_ ), .B1(\RegFile/_3599_ ), .B2(\RegFile/_2177_ ), .C1(\RegFile/_3567_ ), .C2(\RegFile/_2228_ ), .ZN(\RegFile/_2244_ ) );
AOI22_X1 \RegFile/_6321_ ( .A1(\RegFile/_2155_ ), .A2(\RegFile/_3535_ ), .B1(\RegFile/_3311_ ), .B2(\RegFile/_2121_ ), .ZN(\RegFile/_2245_ ) );
AOI22_X1 \RegFile/_6322_ ( .A1(\RegFile/_3343_ ), .A2(\RegFile/_2018_ ), .B1(\RegFile/_2081_ ), .B2(\RegFile/_3375_ ), .ZN(\RegFile/_2246_ ) );
AND3_X1 \RegFile/_6323_ ( .A1(\RegFile/_2040_ ), .A2(\RegFile/_2041_ ), .A3(\RegFile/_3695_ ), .ZN(\RegFile/_2247_ ) );
AOI21_X1 \RegFile/_6324_ ( .A(\RegFile/_2247_ ), .B1(\RegFile/_3727_ ), .B2(\RegFile/_2009_ ), .ZN(\RegFile/_2248_ ) );
AOI22_X1 \RegFile/_6325_ ( .A1(\RegFile/_2085_ ), .A2(\RegFile/_3439_ ), .B1(\RegFile/_3407_ ), .B2(\RegFile/_2086_ ), .ZN(\RegFile/_2249_ ) );
AND4_X1 \RegFile/_6326_ ( .A1(\RegFile/_2245_ ), .A2(\RegFile/_2246_ ), .A3(\RegFile/_2248_ ), .A4(\RegFile/_2249_ ), .ZN(\RegFile/_2250_ ) );
NAND3_X1 \RegFile/_6327_ ( .A1(\RegFile/_2096_ ), .A2(\RegFile/_2161_ ), .A3(\RegFile/_3791_ ), .ZN(\RegFile/_2251_ ) );
NAND3_X1 \RegFile/_6328_ ( .A1(\RegFile/_2096_ ), .A2(\RegFile/_3759_ ), .A3(\RegFile/_2163_ ), .ZN(\RegFile/_2252_ ) );
NAND3_X1 \RegFile/_6329_ ( .A1(\RegFile/_2166_ ), .A2(\RegFile/_2170_ ), .A3(\RegFile/_3503_ ), .ZN(\RegFile/_2253_ ) );
BUF_X4 \RegFile/_6330_ ( .A(\RegFile/_2027_ ), .Z(\RegFile/_2254_ ) );
BUF_X4 \RegFile/_6331_ ( .A(\RegFile/_2028_ ), .Z(\RegFile/_2255_ ) );
NAND3_X1 \RegFile/_6332_ ( .A1(\RegFile/_2254_ ), .A2(\RegFile/_3471_ ), .A3(\RegFile/_2255_ ), .ZN(\RegFile/_2256_ ) );
AND4_X1 \RegFile/_6333_ ( .A1(\RegFile/_2251_ ), .A2(\RegFile/_2252_ ), .A3(\RegFile/_2253_ ), .A4(\RegFile/_2256_ ), .ZN(\RegFile/_2257_ ) );
NAND4_X1 \RegFile/_6334_ ( .A1(\RegFile/_2244_ ), .A2(\RegFile/_2063_ ), .A3(\RegFile/_2250_ ), .A4(\RegFile/_2257_ ), .ZN(\RegFile/_2258_ ) );
OR3_X1 \RegFile/_6335_ ( .A1(\RegFile/_2067_ ), .A2(\RegFile/_2069_ ), .A3(\RegFile/_0745_ ), .ZN(\RegFile/_2259_ ) );
NAND2_X2 \RegFile/_6336_ ( .A1(\RegFile/_2258_ ), .A2(\RegFile/_2259_ ), .ZN(\RegFile/_2260_ ) );
BUF_X4 \RegFile/_6337_ ( .A(\RegFile/_2260_ ), .Z(\RegFile/_2261_ ) );
AOI21_X1 \RegFile/_6338_ ( .A(\RegFile/_2241_ ), .B1(\RegFile/_2261_ ), .B2(\RegFile/_2075_ ), .ZN(\RegFile/_0615_ ) );
NAND2_X1 \RegFile/_6339_ ( .A1(\RegFile/_2077_ ), .A2(\RegFile/_3504_ ), .ZN(\RegFile/_2262_ ) );
NAND3_X1 \RegFile/_6340_ ( .A1(\RegFile/_2034_ ), .A2(\RegFile/_2091_ ), .A3(\RegFile/_3312_ ), .ZN(\RegFile/_2263_ ) );
OAI21_X1 \RegFile/_6341_ ( .A(\RegFile/_2263_ ), .B1(\RegFile/_2182_ ), .B2(\RegFile/_0977_ ), .ZN(\RegFile/_2264_ ) );
AOI221_X1 \RegFile/_6342_ ( .A(\RegFile/_2264_ ), .B1(\RegFile/_3600_ ), .B2(\RegFile/_2177_ ), .C1(\RegFile/_3568_ ), .C2(\RegFile/_2228_ ), .ZN(\RegFile/_2265_ ) );
AOI22_X1 \RegFile/_6343_ ( .A1(\RegFile/_2085_ ), .A2(\RegFile/_3440_ ), .B1(\RegFile/_2053_ ), .B2(\RegFile/_3632_ ), .ZN(\RegFile/_2266_ ) );
AOI22_X1 \RegFile/_6344_ ( .A1(\RegFile/_2048_ ), .A2(\RegFile/_3536_ ), .B1(\RegFile/_3408_ ), .B2(\RegFile/_2086_ ), .ZN(\RegFile/_2267_ ) );
BUF_X4 \RegFile/_6345_ ( .A(\RegFile/_2001_ ), .Z(\RegFile/_2268_ ) );
NAND3_X1 \RegFile/_6346_ ( .A1(\RegFile/_2268_ ), .A2(\RegFile/_3344_ ), .A3(\RegFile/_2254_ ), .ZN(\RegFile/_2269_ ) );
AND4_X1 \RegFile/_6347_ ( .A1(\RegFile/_2062_ ), .A2(\RegFile/_2266_ ), .A3(\RegFile/_2267_ ), .A4(\RegFile/_2269_ ), .ZN(\RegFile/_2270_ ) );
AND3_X1 \RegFile/_6348_ ( .A1(\RegFile/_2220_ ), .A2(\RegFile/_2106_ ), .A3(\RegFile/_3696_ ), .ZN(\RegFile/_2271_ ) );
AOI221_X4 \RegFile/_6349_ ( .A(\RegFile/_2271_ ), .B1(\RegFile/_2008_ ), .B2(\RegFile/_3728_ ), .C1(\RegFile/_3792_ ), .C2(\RegFile/_2014_ ), .ZN(\RegFile/_2272_ ) );
NAND3_X1 \RegFile/_6350_ ( .A1(\RegFile/_2166_ ), .A2(\RegFile/_2170_ ), .A3(\RegFile/_3504_ ), .ZN(\RegFile/_2273_ ) );
NAND3_X1 \RegFile/_6351_ ( .A1(\RegFile/_2268_ ), .A2(\RegFile/_3760_ ), .A3(\RegFile/_2163_ ), .ZN(\RegFile/_2274_ ) );
NAND3_X1 \RegFile/_6352_ ( .A1(\RegFile/_2268_ ), .A2(\RegFile/_3376_ ), .A3(\RegFile/_1989_ ), .ZN(\RegFile/_2275_ ) );
NAND3_X1 \RegFile/_6353_ ( .A1(\RegFile/_2254_ ), .A2(\RegFile/_3472_ ), .A3(\RegFile/_2255_ ), .ZN(\RegFile/_2276_ ) );
AND4_X1 \RegFile/_6354_ ( .A1(\RegFile/_2273_ ), .A2(\RegFile/_2274_ ), .A3(\RegFile/_2275_ ), .A4(\RegFile/_2276_ ), .ZN(\RegFile/_2277_ ) );
NAND4_X2 \RegFile/_6355_ ( .A1(\RegFile/_2265_ ), .A2(\RegFile/_2270_ ), .A3(\RegFile/_2272_ ), .A4(\RegFile/_2277_ ), .ZN(\RegFile/_2278_ ) );
OR3_X1 \RegFile/_6356_ ( .A1(\RegFile/_2067_ ), .A2(\RegFile/_2069_ ), .A3(\RegFile/_0746_ ), .ZN(\RegFile/_2279_ ) );
NAND2_X2 \RegFile/_6357_ ( .A1(\RegFile/_2278_ ), .A2(\RegFile/_2279_ ), .ZN(\RegFile/_2280_ ) );
OAI21_X1 \RegFile/_6358_ ( .A(\RegFile/_2262_ ), .B1(\RegFile/_2280_ ), .B2(\RegFile/_2114_ ), .ZN(\RegFile/_0616_ ) );
NAND2_X1 \RegFile/_6359_ ( .A1(\RegFile/_2077_ ), .A2(\RegFile/_3505_ ), .ZN(\RegFile/_2281_ ) );
INV_X1 \RegFile/_6360_ ( .A(\RegFile/_3665_ ), .ZN(\RegFile/_2282_ ) );
OAI22_X1 \RegFile/_6361_ ( .A1(\RegFile/_2182_ ), .A2(\RegFile/_2282_ ), .B1(\RegFile/_2179_ ), .B2(\RegFile/_1004_ ), .ZN(\RegFile/_2283_ ) );
AOI221_X1 \RegFile/_6362_ ( .A(\RegFile/_2283_ ), .B1(\RegFile/_3601_ ), .B2(\RegFile/_2177_ ), .C1(\RegFile/_3569_ ), .C2(\RegFile/_2050_ ), .ZN(\RegFile/_2284_ ) );
AOI22_X1 \RegFile/_6363_ ( .A1(\RegFile/_2048_ ), .A2(\RegFile/_3537_ ), .B1(\RegFile/_3313_ ), .B2(\RegFile/_2083_ ), .ZN(\RegFile/_2285_ ) );
AOI22_X1 \RegFile/_6364_ ( .A1(\RegFile/_3345_ ), .A2(\RegFile/_2127_ ), .B1(\RegFile/_2126_ ), .B2(\RegFile/_3377_ ), .ZN(\RegFile/_2286_ ) );
AND3_X1 \RegFile/_6365_ ( .A1(\RegFile/_2220_ ), .A2(\RegFile/_2090_ ), .A3(\RegFile/_3697_ ), .ZN(\RegFile/_2287_ ) );
AOI21_X1 \RegFile/_6366_ ( .A(\RegFile/_2287_ ), .B1(\RegFile/_3729_ ), .B2(\RegFile/_2009_ ), .ZN(\RegFile/_2288_ ) );
AOI22_X1 \RegFile/_6367_ ( .A1(\RegFile/_2085_ ), .A2(\RegFile/_3441_ ), .B1(\RegFile/_3409_ ), .B2(\RegFile/_2023_ ), .ZN(\RegFile/_2289_ ) );
AND4_X1 \RegFile/_6368_ ( .A1(\RegFile/_2285_ ), .A2(\RegFile/_2286_ ), .A3(\RegFile/_2288_ ), .A4(\RegFile/_2289_ ), .ZN(\RegFile/_2290_ ) );
NAND3_X1 \RegFile/_6369_ ( .A1(\RegFile/_2096_ ), .A2(\RegFile/_2098_ ), .A3(\RegFile/_3793_ ), .ZN(\RegFile/_2291_ ) );
NAND3_X1 \RegFile/_6370_ ( .A1(\RegFile/_2100_ ), .A2(\RegFile/_3761_ ), .A3(\RegFile/_2101_ ), .ZN(\RegFile/_2292_ ) );
NAND3_X1 \RegFile/_6371_ ( .A1(\RegFile/_1989_ ), .A2(\RegFile/_2255_ ), .A3(\RegFile/_3505_ ), .ZN(\RegFile/_2293_ ) );
NAND3_X1 \RegFile/_6372_ ( .A1(\RegFile/_2107_ ), .A2(\RegFile/_3473_ ), .A3(\RegFile/_2104_ ), .ZN(\RegFile/_2294_ ) );
AND4_X1 \RegFile/_6373_ ( .A1(\RegFile/_2291_ ), .A2(\RegFile/_2292_ ), .A3(\RegFile/_2293_ ), .A4(\RegFile/_2294_ ), .ZN(\RegFile/_2295_ ) );
NAND4_X1 \RegFile/_6374_ ( .A1(\RegFile/_2284_ ), .A2(\RegFile/_2089_ ), .A3(\RegFile/_2290_ ), .A4(\RegFile/_2295_ ), .ZN(\RegFile/_2296_ ) );
OR3_X1 \RegFile/_6375_ ( .A1(\RegFile/_2236_ ), .A2(\RegFile/_2237_ ), .A3(\RegFile/_0747_ ), .ZN(\RegFile/_2297_ ) );
NAND2_X1 \RegFile/_6376_ ( .A1(\RegFile/_2296_ ), .A2(\RegFile/_2297_ ), .ZN(\RegFile/_2298_ ) );
BUF_X4 \RegFile/_6377_ ( .A(\RegFile/_2298_ ), .Z(\RegFile/_2299_ ) );
OAI21_X1 \RegFile/_6378_ ( .A(\RegFile/_2281_ ), .B1(\RegFile/_2299_ ), .B2(\RegFile/_2114_ ), .ZN(\RegFile/_0617_ ) );
AOI21_X1 \RegFile/_6379_ ( .A(\RegFile/_3475_ ), .B1(\RegFile/_1991_ ), .B2(\RegFile/_1997_ ), .ZN(\RegFile/_2300_ ) );
AND3_X1 \RegFile/_6380_ ( .A1(\RegFile/_2040_ ), .A2(\RegFile/_2027_ ), .A3(\RegFile/_3667_ ), .ZN(\RegFile/_2301_ ) );
AOI21_X1 \RegFile/_6381_ ( .A(\RegFile/_2301_ ), .B1(\RegFile/_3699_ ), .B2(\RegFile/_2152_ ), .ZN(\RegFile/_2302_ ) );
AOI22_X1 \RegFile/_6382_ ( .A1(\RegFile/_3315_ ), .A2(\RegFile/_2018_ ), .B1(\RegFile/_2081_ ), .B2(\RegFile/_3347_ ), .ZN(\RegFile/_2303_ ) );
AOI22_X1 \RegFile/_6383_ ( .A1(\RegFile/_2155_ ), .A2(\RegFile/_3507_ ), .B1(\RegFile/_3283_ ), .B2(\RegFile/_2121_ ), .ZN(\RegFile/_2304_ ) );
AOI22_X1 \RegFile/_6384_ ( .A1(\RegFile/_2031_ ), .A2(\RegFile/_3411_ ), .B1(\RegFile/_3379_ ), .B2(\RegFile/_2086_ ), .ZN(\RegFile/_2305_ ) );
AND4_X1 \RegFile/_6385_ ( .A1(\RegFile/_2302_ ), .A2(\RegFile/_2303_ ), .A3(\RegFile/_2304_ ), .A4(\RegFile/_2305_ ), .ZN(\RegFile/_2306_ ) );
NAND3_X1 \RegFile/_6386_ ( .A1(\RegFile/_2041_ ), .A2(\RegFile/_3539_ ), .A3(\RegFile/_2091_ ), .ZN(\RegFile/_2307_ ) );
NAND3_X1 \RegFile/_6387_ ( .A1(\RegFile/_1988_ ), .A2(\RegFile/_2091_ ), .A3(\RegFile/_3571_ ), .ZN(\RegFile/_2308_ ) );
NAND2_X1 \RegFile/_6388_ ( .A1(\RegFile/_2307_ ), .A2(\RegFile/_2308_ ), .ZN(\RegFile/_2309_ ) );
AOI221_X4 \RegFile/_6389_ ( .A(\RegFile/_2309_ ), .B1(\RegFile/_3603_ ), .B2(\RegFile/_2134_ ), .C1(\RegFile/_3635_ ), .C2(\RegFile/_2133_ ), .ZN(\RegFile/_2310_ ) );
NAND3_X1 \RegFile/_6390_ ( .A1(\RegFile/_2041_ ), .A2(\RegFile/_3443_ ), .A3(\RegFile/_2103_ ), .ZN(\RegFile/_2311_ ) );
NAND3_X1 \RegFile/_6391_ ( .A1(\RegFile/_1988_ ), .A2(\RegFile/_1994_ ), .A3(\RegFile/_3475_ ), .ZN(\RegFile/_2312_ ) );
NAND2_X1 \RegFile/_6392_ ( .A1(\RegFile/_2311_ ), .A2(\RegFile/_2312_ ), .ZN(\RegFile/_2313_ ) );
AOI221_X4 \RegFile/_6393_ ( .A(\RegFile/_2313_ ), .B1(\RegFile/_2130_ ), .B2(\RegFile/_3763_ ), .C1(\RegFile/_3731_ ), .C2(\RegFile/_2131_ ), .ZN(\RegFile/_2314_ ) );
NAND4_X1 \RegFile/_6394_ ( .A1(\RegFile/_2306_ ), .A2(\RegFile/_2063_ ), .A3(\RegFile/_2310_ ), .A4(\RegFile/_2314_ ), .ZN(\RegFile/_2315_ ) );
OR3_X1 \RegFile/_6395_ ( .A1(\RegFile/_2067_ ), .A2(\RegFile/_2069_ ), .A3(\RegFile/_0717_ ), .ZN(\RegFile/_2316_ ) );
NAND2_X1 \RegFile/_6396_ ( .A1(\RegFile/_2315_ ), .A2(\RegFile/_2316_ ), .ZN(\RegFile/_2317_ ) );
BUF_X4 \RegFile/_6397_ ( .A(\RegFile/_2317_ ), .Z(\RegFile/_2318_ ) );
AOI21_X1 \RegFile/_6398_ ( .A(\RegFile/_2300_ ), .B1(\RegFile/_2318_ ), .B2(\RegFile/_2075_ ), .ZN(\RegFile/_0618_ ) );
AOI21_X1 \RegFile/_6399_ ( .A(\RegFile/_3476_ ), .B1(\RegFile/_1991_ ), .B2(\RegFile/_1997_ ), .ZN(\RegFile/_2319_ ) );
AOI22_X1 \RegFile/_6400_ ( .A1(\RegFile/_2050_ ), .A2(\RegFile/_3540_ ), .B1(\RegFile/_2177_ ), .B2(\RegFile/_3572_ ), .ZN(\RegFile/_2320_ ) );
OAI221_X1 \RegFile/_6401_ ( .A(\RegFile/_2320_ ), .B1(\RegFile/_1653_ ), .B2(\RegFile/_2179_ ), .C1(\RegFile/_1661_ ), .C2(\RegFile/_2182_ ), .ZN(\RegFile/_2321_ ) );
AOI22_X1 \RegFile/_6402_ ( .A1(\RegFile/_3316_ ), .A2(\RegFile/_2017_ ), .B1(\RegFile/_2126_ ), .B2(\RegFile/_3348_ ), .ZN(\RegFile/_2322_ ) );
AND3_X1 \RegFile/_6403_ ( .A1(\RegFile/_2117_ ), .A2(\RegFile/_2026_ ), .A3(\RegFile/_3668_ ), .ZN(\RegFile/_2323_ ) );
AOI21_X1 \RegFile/_6404_ ( .A(\RegFile/_2323_ ), .B1(\RegFile/_3700_ ), .B2(\RegFile/_2008_ ), .ZN(\RegFile/_2324_ ) );
AOI22_X1 \RegFile/_6405_ ( .A1(\RegFile/_2120_ ), .A2(\RegFile/_3508_ ), .B1(\RegFile/_3284_ ), .B2(\RegFile/_2059_ ), .ZN(\RegFile/_2325_ ) );
AOI22_X1 \RegFile/_6406_ ( .A1(\RegFile/_2188_ ), .A2(\RegFile/_3412_ ), .B1(\RegFile/_3380_ ), .B2(\RegFile/_2023_ ), .ZN(\RegFile/_2326_ ) );
NAND4_X1 \RegFile/_6407_ ( .A1(\RegFile/_2322_ ), .A2(\RegFile/_2324_ ), .A3(\RegFile/_2325_ ), .A4(\RegFile/_2326_ ), .ZN(\RegFile/_2327_ ) );
NAND3_X1 \RegFile/_6408_ ( .A1(\RegFile/_2100_ ), .A2(\RegFile/_2097_ ), .A3(\RegFile/_3764_ ), .ZN(\RegFile/_2328_ ) );
NAND3_X1 \RegFile/_6409_ ( .A1(\RegFile/_2159_ ), .A2(\RegFile/_3732_ ), .A3(\RegFile/_2101_ ), .ZN(\RegFile/_2329_ ) );
NAND3_X1 \RegFile/_6410_ ( .A1(\RegFile/_2165_ ), .A2(\RegFile/_1995_ ), .A3(\RegFile/_3476_ ), .ZN(\RegFile/_2330_ ) );
NAND3_X1 \RegFile/_6411_ ( .A1(\RegFile/_2168_ ), .A2(\RegFile/_3444_ ), .A3(\RegFile/_1995_ ), .ZN(\RegFile/_2331_ ) );
NAND4_X1 \RegFile/_6412_ ( .A1(\RegFile/_2328_ ), .A2(\RegFile/_2329_ ), .A3(\RegFile/_2330_ ), .A4(\RegFile/_2331_ ), .ZN(\RegFile/_2332_ ) );
NOR4_X1 \RegFile/_6413_ ( .A1(\RegFile/_2321_ ), .A2(\RegFile/_2327_ ), .A3(\RegFile/_2061_ ), .A4(\RegFile/_2332_ ), .ZN(\RegFile/_2333_ ) );
AOI211_X4 \RegFile/_6414_ ( .A(\RegFile/_2068_ ), .B(\RegFile/_0718_ ), .C1(\RegFile/_2035_ ), .C2(\RegFile/_2038_ ), .ZN(\RegFile/_2334_ ) );
OR2_X1 \RegFile/_6415_ ( .A1(\RegFile/_2333_ ), .A2(\RegFile/_2334_ ), .ZN(\RegFile/_2335_ ) );
BUF_X4 \RegFile/_6416_ ( .A(\RegFile/_2335_ ), .Z(\RegFile/_2336_ ) );
AOI21_X1 \RegFile/_6417_ ( .A(\RegFile/_2319_ ), .B1(\RegFile/_2336_ ), .B2(\RegFile/_2075_ ), .ZN(\RegFile/_0619_ ) );
AOI21_X1 \RegFile/_6418_ ( .A(\RegFile/_3477_ ), .B1(\RegFile/_1991_ ), .B2(\RegFile/_1997_ ), .ZN(\RegFile/_2337_ ) );
BUF_X4 \RegFile/_6419_ ( .A(\RegFile/_2117_ ), .Z(\RegFile/_2338_ ) );
AND3_X1 \RegFile/_6420_ ( .A1(\RegFile/_2338_ ), .A2(\RegFile/_2168_ ), .A3(\RegFile/_3669_ ), .ZN(\RegFile/_2339_ ) );
AOI21_X1 \RegFile/_6421_ ( .A(\RegFile/_2339_ ), .B1(\RegFile/_3701_ ), .B2(\RegFile/_2152_ ), .ZN(\RegFile/_2340_ ) );
AOI22_X1 \RegFile/_6422_ ( .A1(\RegFile/_3317_ ), .A2(\RegFile/_2206_ ), .B1(\RegFile/_2021_ ), .B2(\RegFile/_3349_ ), .ZN(\RegFile/_2341_ ) );
AOI22_X1 \RegFile/_6423_ ( .A1(\RegFile/_2155_ ), .A2(\RegFile/_3509_ ), .B1(\RegFile/_3285_ ), .B2(\RegFile/_2066_ ), .ZN(\RegFile/_2342_ ) );
AOI22_X1 \RegFile/_6424_ ( .A1(\RegFile/_2031_ ), .A2(\RegFile/_3413_ ), .B1(\RegFile/_3381_ ), .B2(\RegFile/_2024_ ), .ZN(\RegFile/_2343_ ) );
AND4_X1 \RegFile/_6425_ ( .A1(\RegFile/_2340_ ), .A2(\RegFile/_2341_ ), .A3(\RegFile/_2342_ ), .A4(\RegFile/_2343_ ), .ZN(\RegFile/_2344_ ) );
NAND3_X1 \RegFile/_6426_ ( .A1(\RegFile/_2027_ ), .A2(\RegFile/_3541_ ), .A3(\RegFile/_2038_ ), .ZN(\RegFile/_2345_ ) );
NAND3_X1 \RegFile/_6427_ ( .A1(\RegFile/_2165_ ), .A2(\RegFile/_2091_ ), .A3(\RegFile/_3573_ ), .ZN(\RegFile/_2346_ ) );
NAND2_X1 \RegFile/_6428_ ( .A1(\RegFile/_2345_ ), .A2(\RegFile/_2346_ ), .ZN(\RegFile/_2347_ ) );
AOI221_X4 \RegFile/_6429_ ( .A(\RegFile/_2347_ ), .B1(\RegFile/_3605_ ), .B2(\RegFile/_2134_ ), .C1(\RegFile/_3637_ ), .C2(\RegFile/_2045_ ), .ZN(\RegFile/_2348_ ) );
NAND3_X1 \RegFile/_6430_ ( .A1(\RegFile/_2160_ ), .A2(\RegFile/_2161_ ), .A3(\RegFile/_3765_ ), .ZN(\RegFile/_2349_ ) );
NAND3_X1 \RegFile/_6431_ ( .A1(\RegFile/_2160_ ), .A2(\RegFile/_3733_ ), .A3(\RegFile/_2163_ ), .ZN(\RegFile/_2350_ ) );
NAND3_X1 \RegFile/_6432_ ( .A1(\RegFile/_2166_ ), .A2(\RegFile/_1996_ ), .A3(\RegFile/_3477_ ), .ZN(\RegFile/_2351_ ) );
NAND3_X1 \RegFile/_6433_ ( .A1(\RegFile/_2169_ ), .A2(\RegFile/_3445_ ), .A3(\RegFile/_2170_ ), .ZN(\RegFile/_2352_ ) );
AND4_X1 \RegFile/_6434_ ( .A1(\RegFile/_2349_ ), .A2(\RegFile/_2350_ ), .A3(\RegFile/_2351_ ), .A4(\RegFile/_2352_ ), .ZN(\RegFile/_2353_ ) );
NAND4_X1 \RegFile/_6435_ ( .A1(\RegFile/_2344_ ), .A2(\RegFile/_2063_ ), .A3(\RegFile/_2348_ ), .A4(\RegFile/_2353_ ), .ZN(\RegFile/_2354_ ) );
OR3_X2 \RegFile/_6436_ ( .A1(\RegFile/_2067_ ), .A2(\RegFile/_2069_ ), .A3(\RegFile/_0719_ ), .ZN(\RegFile/_2355_ ) );
NAND2_X2 \RegFile/_6437_ ( .A1(\RegFile/_2354_ ), .A2(\RegFile/_2355_ ), .ZN(\RegFile/_2356_ ) );
AOI21_X1 \RegFile/_6438_ ( .A(\RegFile/_2337_ ), .B1(\RegFile/_2356_ ), .B2(\RegFile/_2075_ ), .ZN(\RegFile/_0620_ ) );
BUF_X4 \RegFile/_6439_ ( .A(\RegFile/_1996_ ), .Z(\RegFile/_2357_ ) );
AOI21_X1 \RegFile/_6440_ ( .A(\RegFile/_3478_ ), .B1(\RegFile/_1991_ ), .B2(\RegFile/_2357_ ), .ZN(\RegFile/_2358_ ) );
AOI22_X1 \RegFile/_6441_ ( .A1(\RegFile/_2045_ ), .A2(\RegFile/_3638_ ), .B1(\RegFile/_2053_ ), .B2(\RegFile/_3606_ ), .ZN(\RegFile/_2359_ ) );
INV_X1 \RegFile/_6442_ ( .A(\RegFile/_3574_ ), .ZN(\RegFile/_2360_ ) );
INV_X1 \RegFile/_6443_ ( .A(\RegFile/_3542_ ), .ZN(\RegFile/_2361_ ) );
BUF_X4 \RegFile/_6444_ ( .A(\RegFile/_2144_ ), .Z(\RegFile/_2362_ ) );
OAI221_X1 \RegFile/_6445_ ( .A(\RegFile/_2359_ ), .B1(\RegFile/_2360_ ), .B2(\RegFile/_2146_ ), .C1(\RegFile/_2361_ ), .C2(\RegFile/_2362_ ), .ZN(\RegFile/_2363_ ) );
AOI22_X1 \RegFile/_6446_ ( .A1(\RegFile/_3318_ ), .A2(\RegFile/_2018_ ), .B1(\RegFile/_2081_ ), .B2(\RegFile/_3350_ ), .ZN(\RegFile/_2364_ ) );
AND3_X1 \RegFile/_6447_ ( .A1(\RegFile/_2220_ ), .A2(\RegFile/_2041_ ), .A3(\RegFile/_3670_ ), .ZN(\RegFile/_2365_ ) );
AOI21_X1 \RegFile/_6448_ ( .A(\RegFile/_2365_ ), .B1(\RegFile/_3702_ ), .B2(\RegFile/_2009_ ), .ZN(\RegFile/_2366_ ) );
AOI22_X1 \RegFile/_6449_ ( .A1(\RegFile/_2120_ ), .A2(\RegFile/_3510_ ), .B1(\RegFile/_3286_ ), .B2(\RegFile/_2083_ ), .ZN(\RegFile/_2367_ ) );
AOI22_X1 \RegFile/_6450_ ( .A1(\RegFile/_2188_ ), .A2(\RegFile/_3414_ ), .B1(\RegFile/_3382_ ), .B2(\RegFile/_2023_ ), .ZN(\RegFile/_2368_ ) );
NAND4_X1 \RegFile/_6451_ ( .A1(\RegFile/_2364_ ), .A2(\RegFile/_2366_ ), .A3(\RegFile/_2367_ ), .A4(\RegFile/_2368_ ), .ZN(\RegFile/_2369_ ) );
NAND3_X1 \RegFile/_6452_ ( .A1(\RegFile/_2100_ ), .A2(\RegFile/_2098_ ), .A3(\RegFile/_3766_ ), .ZN(\RegFile/_2370_ ) );
NAND3_X1 \RegFile/_6453_ ( .A1(\RegFile/_2100_ ), .A2(\RegFile/_3734_ ), .A3(\RegFile/_2101_ ), .ZN(\RegFile/_2371_ ) );
NAND3_X1 \RegFile/_6454_ ( .A1(\RegFile/_1989_ ), .A2(\RegFile/_2104_ ), .A3(\RegFile/_3478_ ), .ZN(\RegFile/_2372_ ) );
NAND3_X1 \RegFile/_6455_ ( .A1(\RegFile/_2107_ ), .A2(\RegFile/_3446_ ), .A3(\RegFile/_2104_ ), .ZN(\RegFile/_2373_ ) );
NAND4_X1 \RegFile/_6456_ ( .A1(\RegFile/_2370_ ), .A2(\RegFile/_2371_ ), .A3(\RegFile/_2372_ ), .A4(\RegFile/_2373_ ), .ZN(\RegFile/_2374_ ) );
NOR4_X1 \RegFile/_6457_ ( .A1(\RegFile/_2363_ ), .A2(\RegFile/_2369_ ), .A3(\RegFile/_2061_ ), .A4(\RegFile/_2374_ ), .ZN(\RegFile/_2375_ ) );
BUF_X4 \RegFile/_6458_ ( .A(\RegFile/_2038_ ), .Z(\RegFile/_2376_ ) );
AOI211_X4 \RegFile/_6459_ ( .A(\RegFile/_2068_ ), .B(\RegFile/_0720_ ), .C1(\RegFile/_2035_ ), .C2(\RegFile/_2376_ ), .ZN(\RegFile/_2377_ ) );
OR2_X2 \RegFile/_6460_ ( .A1(\RegFile/_2375_ ), .A2(\RegFile/_2377_ ), .ZN(\RegFile/_2378_ ) );
BUF_X4 \RegFile/_6461_ ( .A(\RegFile/_2378_ ), .Z(\RegFile/_2379_ ) );
AOI21_X1 \RegFile/_6462_ ( .A(\RegFile/_2358_ ), .B1(\RegFile/_2379_ ), .B2(\RegFile/_2075_ ), .ZN(\RegFile/_0621_ ) );
BUF_X4 \RegFile/_6463_ ( .A(\RegFile/_1990_ ), .Z(\RegFile/_2380_ ) );
AOI21_X1 \RegFile/_6464_ ( .A(\RegFile/_3479_ ), .B1(\RegFile/_2380_ ), .B2(\RegFile/_2357_ ), .ZN(\RegFile/_2381_ ) );
NAND3_X1 \RegFile/_6465_ ( .A1(\RegFile/_2338_ ), .A2(\RegFile/_3703_ ), .A3(\RegFile/_1990_ ), .ZN(\RegFile/_2382_ ) );
NAND3_X1 \RegFile/_6466_ ( .A1(\RegFile/_2012_ ), .A2(\RegFile/_3415_ ), .A3(\RegFile/_1993_ ), .ZN(\RegFile/_2383_ ) );
NAND3_X1 \RegFile/_6467_ ( .A1(\RegFile/_1993_ ), .A2(\RegFile/_2003_ ), .A3(\RegFile/_3383_ ), .ZN(\RegFile/_2384_ ) );
NAND2_X1 \RegFile/_6468_ ( .A1(\RegFile/_2383_ ), .A2(\RegFile/_2384_ ), .ZN(\RegFile/_2385_ ) );
AOI221_X4 \RegFile/_6469_ ( .A(\RegFile/_2385_ ), .B1(\RegFile/_3351_ ), .B2(\RegFile/_2020_ ), .C1(\RegFile/_3319_ ), .C2(\RegFile/_2017_ ), .ZN(\RegFile/_2386_ ) );
NAND3_X1 \RegFile/_6470_ ( .A1(\RegFile/_2338_ ), .A2(\RegFile/_2169_ ), .A3(\RegFile/_3671_ ), .ZN(\RegFile/_2387_ ) );
AOI22_X1 \RegFile/_6471_ ( .A1(\RegFile/_2155_ ), .A2(\RegFile/_3511_ ), .B1(\RegFile/_3287_ ), .B2(\RegFile/_2066_ ), .ZN(\RegFile/_2388_ ) );
AND4_X1 \RegFile/_6472_ ( .A1(\RegFile/_2382_ ), .A2(\RegFile/_2386_ ), .A3(\RegFile/_2387_ ), .A4(\RegFile/_2388_ ), .ZN(\RegFile/_2389_ ) );
INV_X1 \RegFile/_6473_ ( .A(\RegFile/_3575_ ), .ZN(\RegFile/_2390_ ) );
OAI22_X1 \RegFile/_6474_ ( .A1(\RegFile/_2144_ ), .A2(\RegFile/_1701_ ), .B1(\RegFile/_2146_ ), .B2(\RegFile/_2390_ ), .ZN(\RegFile/_2391_ ) );
AOI221_X4 \RegFile/_6475_ ( .A(\RegFile/_2391_ ), .B1(\RegFile/_3639_ ), .B2(\RegFile/_2133_ ), .C1(\RegFile/_3607_ ), .C2(\RegFile/_2053_ ), .ZN(\RegFile/_2392_ ) );
NAND3_X1 \RegFile/_6476_ ( .A1(\RegFile/_2027_ ), .A2(\RegFile/_3447_ ), .A3(\RegFile/_2028_ ), .ZN(\RegFile/_2393_ ) );
NAND3_X1 \RegFile/_6477_ ( .A1(\RegFile/_2165_ ), .A2(\RegFile/_2028_ ), .A3(\RegFile/_3479_ ), .ZN(\RegFile/_2394_ ) );
NAND2_X1 \RegFile/_6478_ ( .A1(\RegFile/_2393_ ), .A2(\RegFile/_2394_ ), .ZN(\RegFile/_2395_ ) );
AOI221_X4 \RegFile/_6479_ ( .A(\RegFile/_2395_ ), .B1(\RegFile/_2130_ ), .B2(\RegFile/_3767_ ), .C1(\RegFile/_3735_ ), .C2(\RegFile/_2005_ ), .ZN(\RegFile/_2396_ ) );
NAND4_X4 \RegFile/_6480_ ( .A1(\RegFile/_2389_ ), .A2(\RegFile/_2063_ ), .A3(\RegFile/_2392_ ), .A4(\RegFile/_2396_ ), .ZN(\RegFile/_2397_ ) );
OR3_X2 \RegFile/_6481_ ( .A1(\RegFile/_2067_ ), .A2(\RegFile/_2069_ ), .A3(\RegFile/_0721_ ), .ZN(\RegFile/_2398_ ) );
NAND2_X2 \RegFile/_6482_ ( .A1(\RegFile/_2397_ ), .A2(\RegFile/_2398_ ), .ZN(\RegFile/_2399_ ) );
BUF_X4 \RegFile/_6483_ ( .A(\RegFile/_2074_ ), .Z(\RegFile/_2400_ ) );
AOI21_X1 \RegFile/_6484_ ( .A(\RegFile/_2381_ ), .B1(\RegFile/_2399_ ), .B2(\RegFile/_2400_ ), .ZN(\RegFile/_0622_ ) );
AOI21_X1 \RegFile/_6485_ ( .A(\RegFile/_3480_ ), .B1(\RegFile/_2380_ ), .B2(\RegFile/_2357_ ), .ZN(\RegFile/_2401_ ) );
AOI22_X1 \RegFile/_6486_ ( .A1(\RegFile/_3320_ ), .A2(\RegFile/_2017_ ), .B1(\RegFile/_2020_ ), .B2(\RegFile/_3352_ ), .ZN(\RegFile/_2402_ ) );
NAND3_X1 \RegFile/_6487_ ( .A1(\RegFile/_1995_ ), .A2(\RegFile/_2101_ ), .A3(\RegFile/_3384_ ), .ZN(\RegFile/_2403_ ) );
INV_X2 \RegFile/_6488_ ( .A(\RegFile/_2188_ ), .ZN(\RegFile/_2404_ ) );
OAI211_X2 \RegFile/_6489_ ( .A(\RegFile/_2402_ ), .B(\RegFile/_2403_ ), .C1(\RegFile/_1097_ ), .C2(\RegFile/_2404_ ), .ZN(\RegFile/_2405_ ) );
AOI22_X1 \RegFile/_6490_ ( .A1(\RegFile/_3768_ ), .A2(\RegFile/_2130_ ), .B1(\RegFile/_2004_ ), .B2(\RegFile/_3736_ ), .ZN(\RegFile/_2406_ ) );
AOI22_X1 \RegFile/_6491_ ( .A1(\RegFile/_2050_ ), .A2(\RegFile/_3544_ ), .B1(\RegFile/_2177_ ), .B2(\RegFile/_3576_ ), .ZN(\RegFile/_2407_ ) );
AOI22_X1 \RegFile/_6492_ ( .A1(\RegFile/_2044_ ), .A2(\RegFile/_3640_ ), .B1(\RegFile/_2134_ ), .B2(\RegFile/_3608_ ), .ZN(\RegFile/_2408_ ) );
AND3_X1 \RegFile/_6493_ ( .A1(\RegFile/_2026_ ), .A2(\RegFile/_3448_ ), .A3(\RegFile/_1994_ ), .ZN(\RegFile/_2409_ ) );
AOI21_X1 \RegFile/_6494_ ( .A(\RegFile/_2409_ ), .B1(\RegFile/_3480_ ), .B2(\RegFile/_2074_ ), .ZN(\RegFile/_2410_ ) );
NAND4_X1 \RegFile/_6495_ ( .A1(\RegFile/_2406_ ), .A2(\RegFile/_2407_ ), .A3(\RegFile/_2408_ ), .A4(\RegFile/_2410_ ), .ZN(\RegFile/_2411_ ) );
AND3_X1 \RegFile/_6496_ ( .A1(\RegFile/_2003_ ), .A2(\RegFile/_2037_ ), .A3(\RegFile/_3288_ ), .ZN(\RegFile/_2412_ ) );
AND3_X1 \RegFile/_6497_ ( .A1(\RegFile/_2012_ ), .A2(\RegFile/_3512_ ), .A3(\RegFile/_2037_ ), .ZN(\RegFile/_2413_ ) );
AND3_X1 \RegFile/_6498_ ( .A1(\RegFile/_2006_ ), .A2(\RegFile/_2026_ ), .A3(\RegFile/_3672_ ), .ZN(\RegFile/_2414_ ) );
AND3_X4 \RegFile/_6499_ ( .A1(\RegFile/_2006_ ), .A2(\RegFile/_3704_ ), .A3(\RegFile/_1988_ ), .ZN(\RegFile/_2415_ ) );
OR4_X4 \RegFile/_6500_ ( .A1(\RegFile/_2412_ ), .A2(\RegFile/_2413_ ), .A3(\RegFile/_2414_ ), .A4(\RegFile/_2415_ ), .ZN(\RegFile/_2416_ ) );
OR4_X4 \RegFile/_6501_ ( .A1(\RegFile/_2061_ ), .A2(\RegFile/_2405_ ), .A3(\RegFile/_2411_ ), .A4(\RegFile/_2416_ ), .ZN(\RegFile/_2417_ ) );
OR3_X1 \RegFile/_6502_ ( .A1(\RegFile/_2236_ ), .A2(\RegFile/_2237_ ), .A3(\RegFile/_0722_ ), .ZN(\RegFile/_2418_ ) );
NAND2_X4 \RegFile/_6503_ ( .A1(\RegFile/_2417_ ), .A2(\RegFile/_2418_ ), .ZN(\RegFile/_2419_ ) );
BUF_X8 \RegFile/_6504_ ( .A(\RegFile/_2419_ ), .Z(\RegFile/_2420_ ) );
AOI21_X1 \RegFile/_6505_ ( .A(\RegFile/_2401_ ), .B1(\RegFile/_2420_ ), .B2(\RegFile/_2400_ ), .ZN(\RegFile/_0623_ ) );
AOI21_X1 \RegFile/_6506_ ( .A(\RegFile/_3481_ ), .B1(\RegFile/_2380_ ), .B2(\RegFile/_2357_ ), .ZN(\RegFile/_2421_ ) );
AND3_X1 \RegFile/_6507_ ( .A1(\RegFile/_2040_ ), .A2(\RegFile/_2027_ ), .A3(\RegFile/_3673_ ), .ZN(\RegFile/_2422_ ) );
AOI21_X1 \RegFile/_6508_ ( .A(\RegFile/_2422_ ), .B1(\RegFile/_3705_ ), .B2(\RegFile/_2009_ ), .ZN(\RegFile/_2423_ ) );
AOI22_X1 \RegFile/_6509_ ( .A1(\RegFile/_3321_ ), .A2(\RegFile/_2018_ ), .B1(\RegFile/_2081_ ), .B2(\RegFile/_3353_ ), .ZN(\RegFile/_2424_ ) );
AOI22_X1 \RegFile/_6510_ ( .A1(\RegFile/_2048_ ), .A2(\RegFile/_3513_ ), .B1(\RegFile/_3289_ ), .B2(\RegFile/_2083_ ), .ZN(\RegFile/_2425_ ) );
AOI22_X1 \RegFile/_6511_ ( .A1(\RegFile/_2085_ ), .A2(\RegFile/_3417_ ), .B1(\RegFile/_3385_ ), .B2(\RegFile/_2086_ ), .ZN(\RegFile/_2426_ ) );
AND4_X1 \RegFile/_6512_ ( .A1(\RegFile/_2423_ ), .A2(\RegFile/_2424_ ), .A3(\RegFile/_2425_ ), .A4(\RegFile/_2426_ ), .ZN(\RegFile/_2427_ ) );
NAND3_X1 \RegFile/_6513_ ( .A1(\RegFile/_2097_ ), .A2(\RegFile/_3641_ ), .A3(\RegFile/_2117_ ), .ZN(\RegFile/_2428_ ) );
NAND3_X1 \RegFile/_6514_ ( .A1(\RegFile/_2220_ ), .A2(\RegFile/_3609_ ), .A3(\RegFile/_2034_ ), .ZN(\RegFile/_2429_ ) );
NAND2_X1 \RegFile/_6515_ ( .A1(\RegFile/_2428_ ), .A2(\RegFile/_2429_ ), .ZN(\RegFile/_2430_ ) );
AOI221_X4 \RegFile/_6516_ ( .A(\RegFile/_2430_ ), .B1(\RegFile/_3577_ ), .B2(\RegFile/_2177_ ), .C1(\RegFile/_3545_ ), .C2(\RegFile/_2050_ ), .ZN(\RegFile/_2431_ ) );
NAND3_X1 \RegFile/_6517_ ( .A1(\RegFile/_2096_ ), .A2(\RegFile/_2098_ ), .A3(\RegFile/_3769_ ), .ZN(\RegFile/_2432_ ) );
NAND3_X1 \RegFile/_6518_ ( .A1(\RegFile/_2268_ ), .A2(\RegFile/_3737_ ), .A3(\RegFile/_2101_ ), .ZN(\RegFile/_2433_ ) );
NAND3_X1 \RegFile/_6519_ ( .A1(\RegFile/_2166_ ), .A2(\RegFile/_2255_ ), .A3(\RegFile/_3481_ ), .ZN(\RegFile/_2434_ ) );
NAND3_X1 \RegFile/_6520_ ( .A1(\RegFile/_2254_ ), .A2(\RegFile/_3449_ ), .A3(\RegFile/_2255_ ), .ZN(\RegFile/_2435_ ) );
AND4_X1 \RegFile/_6521_ ( .A1(\RegFile/_2432_ ), .A2(\RegFile/_2433_ ), .A3(\RegFile/_2434_ ), .A4(\RegFile/_2435_ ), .ZN(\RegFile/_2436_ ) );
NAND4_X1 \RegFile/_6522_ ( .A1(\RegFile/_2427_ ), .A2(\RegFile/_2089_ ), .A3(\RegFile/_2431_ ), .A4(\RegFile/_2436_ ), .ZN(\RegFile/_2437_ ) );
OR3_X1 \RegFile/_6523_ ( .A1(\RegFile/_2236_ ), .A2(\RegFile/_2237_ ), .A3(\RegFile/_0723_ ), .ZN(\RegFile/_2438_ ) );
NAND2_X1 \RegFile/_6524_ ( .A1(\RegFile/_2437_ ), .A2(\RegFile/_2438_ ), .ZN(\RegFile/_2439_ ) );
BUF_X4 \RegFile/_6525_ ( .A(\RegFile/_2439_ ), .Z(\RegFile/_2440_ ) );
AOI21_X1 \RegFile/_6526_ ( .A(\RegFile/_2421_ ), .B1(\RegFile/_2440_ ), .B2(\RegFile/_2400_ ), .ZN(\RegFile/_0624_ ) );
AOI21_X1 \RegFile/_6527_ ( .A(\RegFile/_3482_ ), .B1(\RegFile/_2380_ ), .B2(\RegFile/_2357_ ), .ZN(\RegFile/_2441_ ) );
AOI22_X1 \RegFile/_6528_ ( .A1(\RegFile/_3770_ ), .A2(\RegFile/_2130_ ), .B1(\RegFile/_2131_ ), .B2(\RegFile/_3738_ ), .ZN(\RegFile/_2442_ ) );
AOI22_X1 \RegFile/_6529_ ( .A1(\RegFile/_2050_ ), .A2(\RegFile/_3546_ ), .B1(\RegFile/_2177_ ), .B2(\RegFile/_3578_ ), .ZN(\RegFile/_2443_ ) );
AOI22_X1 \RegFile/_6530_ ( .A1(\RegFile/_2133_ ), .A2(\RegFile/_3642_ ), .B1(\RegFile/_2134_ ), .B2(\RegFile/_3610_ ), .ZN(\RegFile/_2444_ ) );
AND3_X1 \RegFile/_6531_ ( .A1(\RegFile/_2106_ ), .A2(\RegFile/_3450_ ), .A3(\RegFile/_1994_ ), .ZN(\RegFile/_2445_ ) );
AOI21_X1 \RegFile/_6532_ ( .A(\RegFile/_2445_ ), .B1(\RegFile/_3482_ ), .B2(\RegFile/_2074_ ), .ZN(\RegFile/_2446_ ) );
NAND4_X1 \RegFile/_6533_ ( .A1(\RegFile/_2442_ ), .A2(\RegFile/_2443_ ), .A3(\RegFile/_2444_ ), .A4(\RegFile/_2446_ ), .ZN(\RegFile/_2447_ ) );
AOI22_X1 \RegFile/_6534_ ( .A1(\RegFile/_2120_ ), .A2(\RegFile/_3514_ ), .B1(\RegFile/_3290_ ), .B2(\RegFile/_2059_ ), .ZN(\RegFile/_2448_ ) );
NAND3_X1 \RegFile/_6535_ ( .A1(\RegFile/_2338_ ), .A2(\RegFile/_2107_ ), .A3(\RegFile/_3674_ ), .ZN(\RegFile/_2449_ ) );
OAI211_X2 \RegFile/_6536_ ( .A(\RegFile/_2448_ ), .B(\RegFile/_2449_ ), .C1(\RegFile/_1141_ ), .C2(\RegFile/_2116_ ), .ZN(\RegFile/_2450_ ) );
NAND3_X1 \RegFile/_6537_ ( .A1(\RegFile/_2098_ ), .A2(\RegFile/_3418_ ), .A3(\RegFile/_1995_ ), .ZN(\RegFile/_2451_ ) );
NAND3_X1 \RegFile/_6538_ ( .A1(\RegFile/_2159_ ), .A2(\RegFile/_3354_ ), .A3(\RegFile/_2165_ ), .ZN(\RegFile/_2452_ ) );
NAND3_X1 \RegFile/_6539_ ( .A1(\RegFile/_2159_ ), .A2(\RegFile/_3322_ ), .A3(\RegFile/_2168_ ), .ZN(\RegFile/_2453_ ) );
NAND3_X1 \RegFile/_6540_ ( .A1(\RegFile/_1995_ ), .A2(\RegFile/_2034_ ), .A3(\RegFile/_3386_ ), .ZN(\RegFile/_2454_ ) );
NAND4_X1 \RegFile/_6541_ ( .A1(\RegFile/_2451_ ), .A2(\RegFile/_2452_ ), .A3(\RegFile/_2453_ ), .A4(\RegFile/_2454_ ), .ZN(\RegFile/_2455_ ) );
NOR4_X1 \RegFile/_6542_ ( .A1(\RegFile/_2447_ ), .A2(\RegFile/_2450_ ), .A3(\RegFile/_2061_ ), .A4(\RegFile/_2455_ ), .ZN(\RegFile/_2456_ ) );
AOI211_X4 \RegFile/_6543_ ( .A(\RegFile/_2060_ ), .B(\RegFile/_0724_ ), .C1(\RegFile/_2035_ ), .C2(\RegFile/_2038_ ), .ZN(\RegFile/_2457_ ) );
OR2_X1 \RegFile/_6544_ ( .A1(\RegFile/_2456_ ), .A2(\RegFile/_2457_ ), .ZN(\RegFile/_2458_ ) );
BUF_X4 \RegFile/_6545_ ( .A(\RegFile/_2458_ ), .Z(\RegFile/_2459_ ) );
AOI21_X1 \RegFile/_6546_ ( .A(\RegFile/_2441_ ), .B1(\RegFile/_2459_ ), .B2(\RegFile/_2400_ ), .ZN(\RegFile/_0625_ ) );
NAND2_X1 \RegFile/_6547_ ( .A1(\RegFile/_2077_ ), .A2(\RegFile/_3483_ ), .ZN(\RegFile/_2460_ ) );
OAI22_X1 \RegFile/_6548_ ( .A1(\RegFile/_2116_ ), .A2(\RegFile/_1158_ ), .B1(\RegFile/_2118_ ), .B2(\RegFile/_1155_ ), .ZN(\RegFile/_2461_ ) );
AOI221_X4 \RegFile/_6549_ ( .A(\RegFile/_2461_ ), .B1(\RegFile/_3515_ ), .B2(\RegFile/_2120_ ), .C1(\RegFile/_3291_ ), .C2(\RegFile/_2121_ ), .ZN(\RegFile/_2462_ ) );
NAND3_X1 \RegFile/_6550_ ( .A1(\RegFile/_2001_ ), .A2(\RegFile/_3355_ ), .A3(\RegFile/_1988_ ), .ZN(\RegFile/_2463_ ) );
NAND3_X1 \RegFile/_6551_ ( .A1(\RegFile/_2001_ ), .A2(\RegFile/_3323_ ), .A3(\RegFile/_2106_ ), .ZN(\RegFile/_2464_ ) );
NAND2_X1 \RegFile/_6552_ ( .A1(\RegFile/_2463_ ), .A2(\RegFile/_2464_ ), .ZN(\RegFile/_2465_ ) );
AOI221_X4 \RegFile/_6553_ ( .A(\RegFile/_2465_ ), .B1(\RegFile/_3419_ ), .B2(\RegFile/_2188_ ), .C1(\RegFile/_3387_ ), .C2(\RegFile/_2024_ ), .ZN(\RegFile/_2466_ ) );
AOI22_X1 \RegFile/_6554_ ( .A1(\RegFile/_2050_ ), .A2(\RegFile/_3547_ ), .B1(\RegFile/_2055_ ), .B2(\RegFile/_3579_ ), .ZN(\RegFile/_2467_ ) );
AOI22_X1 \RegFile/_6555_ ( .A1(\RegFile/_3771_ ), .A2(\RegFile/_2130_ ), .B1(\RegFile/_2131_ ), .B2(\RegFile/_3739_ ), .ZN(\RegFile/_2468_ ) );
AOI22_X1 \RegFile/_6556_ ( .A1(\RegFile/_2133_ ), .A2(\RegFile/_3643_ ), .B1(\RegFile/_2134_ ), .B2(\RegFile/_3611_ ), .ZN(\RegFile/_2469_ ) );
AND3_X1 \RegFile/_6557_ ( .A1(\RegFile/_2090_ ), .A2(\RegFile/_3451_ ), .A3(\RegFile/_1994_ ), .ZN(\RegFile/_2470_ ) );
AOI21_X1 \RegFile/_6558_ ( .A(\RegFile/_2470_ ), .B1(\RegFile/_3483_ ), .B2(\RegFile/_2074_ ), .ZN(\RegFile/_2471_ ) );
AND4_X1 \RegFile/_6559_ ( .A1(\RegFile/_2467_ ), .A2(\RegFile/_2468_ ), .A3(\RegFile/_2469_ ), .A4(\RegFile/_2471_ ), .ZN(\RegFile/_2472_ ) );
NAND4_X4 \RegFile/_6560_ ( .A1(\RegFile/_2462_ ), .A2(\RegFile/_2089_ ), .A3(\RegFile/_2466_ ), .A4(\RegFile/_2472_ ), .ZN(\RegFile/_2473_ ) );
OR3_X1 \RegFile/_6561_ ( .A1(\RegFile/_2236_ ), .A2(\RegFile/_2237_ ), .A3(\RegFile/_0725_ ), .ZN(\RegFile/_2474_ ) );
NAND2_X1 \RegFile/_6562_ ( .A1(\RegFile/_2473_ ), .A2(\RegFile/_2474_ ), .ZN(\RegFile/_2475_ ) );
BUF_X4 \RegFile/_6563_ ( .A(\RegFile/_2475_ ), .Z(\RegFile/_2476_ ) );
OAI21_X1 \RegFile/_6564_ ( .A(\RegFile/_2460_ ), .B1(\RegFile/_2476_ ), .B2(\RegFile/_2114_ ), .ZN(\RegFile/_0626_ ) );
NAND2_X1 \RegFile/_6565_ ( .A1(\RegFile/_2077_ ), .A2(\RegFile/_3484_ ), .ZN(\RegFile/_2477_ ) );
AOI22_X1 \RegFile/_6566_ ( .A1(\RegFile/_3324_ ), .A2(\RegFile/_2127_ ), .B1(\RegFile/_2126_ ), .B2(\RegFile/_3356_ ), .ZN(\RegFile/_2478_ ) );
AND3_X1 \RegFile/_6567_ ( .A1(\RegFile/_2117_ ), .A2(\RegFile/_2106_ ), .A3(\RegFile/_3676_ ), .ZN(\RegFile/_2479_ ) );
AOI21_X1 \RegFile/_6568_ ( .A(\RegFile/_2479_ ), .B1(\RegFile/_3708_ ), .B2(\RegFile/_2008_ ), .ZN(\RegFile/_2480_ ) );
AOI22_X1 \RegFile/_6569_ ( .A1(\RegFile/_2120_ ), .A2(\RegFile/_3516_ ), .B1(\RegFile/_3292_ ), .B2(\RegFile/_2083_ ), .ZN(\RegFile/_2481_ ) );
AOI22_X1 \RegFile/_6570_ ( .A1(\RegFile/_2188_ ), .A2(\RegFile/_3420_ ), .B1(\RegFile/_3388_ ), .B2(\RegFile/_2023_ ), .ZN(\RegFile/_2482_ ) );
NAND4_X1 \RegFile/_6571_ ( .A1(\RegFile/_2478_ ), .A2(\RegFile/_2480_ ), .A3(\RegFile/_2481_ ), .A4(\RegFile/_2482_ ), .ZN(\RegFile/_2483_ ) );
AOI22_X1 \RegFile/_6572_ ( .A1(\RegFile/_2044_ ), .A2(\RegFile/_3644_ ), .B1(\RegFile/_2052_ ), .B2(\RegFile/_3612_ ), .ZN(\RegFile/_2484_ ) );
NAND3_X1 \RegFile/_6573_ ( .A1(\RegFile/_2168_ ), .A2(\RegFile/_3548_ ), .A3(\RegFile/_2038_ ), .ZN(\RegFile/_2485_ ) );
OAI211_X2 \RegFile/_6574_ ( .A(\RegFile/_2484_ ), .B(\RegFile/_2485_ ), .C1(\RegFile/_1174_ ), .C2(\RegFile/_2146_ ), .ZN(\RegFile/_2486_ ) );
NAND3_X1 \RegFile/_6575_ ( .A1(\RegFile/_2159_ ), .A2(\RegFile/_2097_ ), .A3(\RegFile/_3772_ ), .ZN(\RegFile/_2487_ ) );
NAND3_X1 \RegFile/_6576_ ( .A1(\RegFile/_2159_ ), .A2(\RegFile/_3740_ ), .A3(\RegFile/_2034_ ), .ZN(\RegFile/_2488_ ) );
NAND3_X1 \RegFile/_6577_ ( .A1(\RegFile/_2165_ ), .A2(\RegFile/_1995_ ), .A3(\RegFile/_3484_ ), .ZN(\RegFile/_2489_ ) );
NAND3_X1 \RegFile/_6578_ ( .A1(\RegFile/_2168_ ), .A2(\RegFile/_3452_ ), .A3(\RegFile/_2028_ ), .ZN(\RegFile/_2490_ ) );
NAND4_X1 \RegFile/_6579_ ( .A1(\RegFile/_2487_ ), .A2(\RegFile/_2488_ ), .A3(\RegFile/_2489_ ), .A4(\RegFile/_2490_ ), .ZN(\RegFile/_2491_ ) );
NOR4_X1 \RegFile/_6580_ ( .A1(\RegFile/_2483_ ), .A2(\RegFile/_2486_ ), .A3(\RegFile/_2061_ ), .A4(\RegFile/_2491_ ), .ZN(\RegFile/_2492_ ) );
AOI211_X4 \RegFile/_6581_ ( .A(\RegFile/_2060_ ), .B(\RegFile/_0726_ ), .C1(\RegFile/_2163_ ), .C2(\RegFile/_2038_ ), .ZN(\RegFile/_2493_ ) );
OR2_X2 \RegFile/_6582_ ( .A1(\RegFile/_2492_ ), .A2(\RegFile/_2493_ ), .ZN(\RegFile/_2494_ ) );
BUF_X4 \RegFile/_6583_ ( .A(\RegFile/_2494_ ), .Z(\RegFile/_2495_ ) );
OAI21_X1 \RegFile/_6584_ ( .A(\RegFile/_2477_ ), .B1(\RegFile/_2495_ ), .B2(\RegFile/_2114_ ), .ZN(\RegFile/_0627_ ) );
AOI21_X1 \RegFile/_6585_ ( .A(\RegFile/_3486_ ), .B1(\RegFile/_2380_ ), .B2(\RegFile/_2357_ ), .ZN(\RegFile/_2496_ ) );
AOI22_X1 \RegFile/_6586_ ( .A1(\RegFile/_3326_ ), .A2(\RegFile/_2127_ ), .B1(\RegFile/_2126_ ), .B2(\RegFile/_3358_ ), .ZN(\RegFile/_2497_ ) );
AND3_X1 \RegFile/_6587_ ( .A1(\RegFile/_2117_ ), .A2(\RegFile/_2026_ ), .A3(\RegFile/_3678_ ), .ZN(\RegFile/_2498_ ) );
AOI21_X1 \RegFile/_6588_ ( .A(\RegFile/_2498_ ), .B1(\RegFile/_3710_ ), .B2(\RegFile/_2008_ ), .ZN(\RegFile/_2499_ ) );
AOI22_X1 \RegFile/_6589_ ( .A1(\RegFile/_2120_ ), .A2(\RegFile/_3518_ ), .B1(\RegFile/_3294_ ), .B2(\RegFile/_2083_ ), .ZN(\RegFile/_2500_ ) );
AOI22_X1 \RegFile/_6590_ ( .A1(\RegFile/_2188_ ), .A2(\RegFile/_3422_ ), .B1(\RegFile/_3390_ ), .B2(\RegFile/_2023_ ), .ZN(\RegFile/_2501_ ) );
NAND4_X1 \RegFile/_6591_ ( .A1(\RegFile/_2497_ ), .A2(\RegFile/_2499_ ), .A3(\RegFile/_2500_ ), .A4(\RegFile/_2501_ ), .ZN(\RegFile/_2502_ ) );
AOI22_X2 \RegFile/_6592_ ( .A1(\RegFile/_2050_ ), .A2(\RegFile/_3550_ ), .B1(\RegFile/_2177_ ), .B2(\RegFile/_3582_ ), .ZN(\RegFile/_2503_ ) );
NAND3_X1 \RegFile/_6593_ ( .A1(\RegFile/_2097_ ), .A2(\RegFile/_3646_ ), .A3(\RegFile/_2338_ ), .ZN(\RegFile/_2504_ ) );
OAI211_X2 \RegFile/_6594_ ( .A(\RegFile/_2503_ ), .B(\RegFile/_2504_ ), .C1(\RegFile/_1806_ ), .C2(\RegFile/_2179_ ), .ZN(\RegFile/_2505_ ) );
NAND3_X1 \RegFile/_6595_ ( .A1(\RegFile/_2159_ ), .A2(\RegFile/_2097_ ), .A3(\RegFile/_3774_ ), .ZN(\RegFile/_2506_ ) );
NAND3_X1 \RegFile/_6596_ ( .A1(\RegFile/_2159_ ), .A2(\RegFile/_3742_ ), .A3(\RegFile/_2034_ ), .ZN(\RegFile/_2507_ ) );
NAND3_X1 \RegFile/_6597_ ( .A1(\RegFile/_2165_ ), .A2(\RegFile/_2028_ ), .A3(\RegFile/_3486_ ), .ZN(\RegFile/_2508_ ) );
NAND3_X1 \RegFile/_6598_ ( .A1(\RegFile/_2168_ ), .A2(\RegFile/_3454_ ), .A3(\RegFile/_2028_ ), .ZN(\RegFile/_2509_ ) );
NAND4_X1 \RegFile/_6599_ ( .A1(\RegFile/_2506_ ), .A2(\RegFile/_2507_ ), .A3(\RegFile/_2508_ ), .A4(\RegFile/_2509_ ), .ZN(\RegFile/_2510_ ) );
NOR4_X2 \RegFile/_6600_ ( .A1(\RegFile/_2502_ ), .A2(\RegFile/_2505_ ), .A3(\RegFile/_2061_ ), .A4(\RegFile/_2510_ ), .ZN(\RegFile/_2511_ ) );
AOI211_X4 \RegFile/_6601_ ( .A(\RegFile/_2060_ ), .B(\RegFile/_0728_ ), .C1(\RegFile/_2163_ ), .C2(\RegFile/_2038_ ), .ZN(\RegFile/_2512_ ) );
OR2_X2 \RegFile/_6602_ ( .A1(\RegFile/_2511_ ), .A2(\RegFile/_2512_ ), .ZN(\RegFile/_2513_ ) );
BUF_X4 \RegFile/_6603_ ( .A(\RegFile/_2513_ ), .Z(\RegFile/_2514_ ) );
AOI21_X1 \RegFile/_6604_ ( .A(\RegFile/_2496_ ), .B1(\RegFile/_2514_ ), .B2(\RegFile/_2400_ ), .ZN(\RegFile/_0628_ ) );
AOI21_X1 \RegFile/_6605_ ( .A(\RegFile/_3487_ ), .B1(\RegFile/_2380_ ), .B2(\RegFile/_2357_ ), .ZN(\RegFile/_2515_ ) );
NAND3_X1 \RegFile/_6606_ ( .A1(\RegFile/_2166_ ), .A2(\RegFile/_2170_ ), .A3(\RegFile/_3487_ ), .ZN(\RegFile/_2516_ ) );
INV_X1 \RegFile/_6607_ ( .A(\RegFile/_3583_ ), .ZN(\RegFile/_2517_ ) );
OAI22_X1 \RegFile/_6608_ ( .A1(\RegFile/_2144_ ), .A2(\RegFile/_1816_ ), .B1(\RegFile/_2145_ ), .B2(\RegFile/_2517_ ), .ZN(\RegFile/_2518_ ) );
AOI221_X1 \RegFile/_6609_ ( .A(\RegFile/_2518_ ), .B1(\RegFile/_3647_ ), .B2(\RegFile/_2044_ ), .C1(\RegFile/_3615_ ), .C2(\RegFile/_2052_ ), .ZN(\RegFile/_2519_ ) );
NAND3_X1 \RegFile/_6610_ ( .A1(\RegFile/_2254_ ), .A2(\RegFile/_3455_ ), .A3(\RegFile/_2170_ ), .ZN(\RegFile/_2520_ ) );
AOI22_X1 \RegFile/_6611_ ( .A1(\RegFile/_3775_ ), .A2(\RegFile/_2014_ ), .B1(\RegFile/_2131_ ), .B2(\RegFile/_3743_ ), .ZN(\RegFile/_2521_ ) );
AND4_X1 \RegFile/_6612_ ( .A1(\RegFile/_2516_ ), .A2(\RegFile/_2519_ ), .A3(\RegFile/_2520_ ), .A4(\RegFile/_2521_ ), .ZN(\RegFile/_2522_ ) );
NAND3_X1 \RegFile/_6613_ ( .A1(\RegFile/_2117_ ), .A2(\RegFile/_2106_ ), .A3(\RegFile/_3679_ ), .ZN(\RegFile/_2523_ ) );
OAI21_X1 \RegFile/_6614_ ( .A(\RegFile/_2523_ ), .B1(\RegFile/_2116_ ), .B2(\RegFile/_1819_ ), .ZN(\RegFile/_2524_ ) );
AOI221_X4 \RegFile/_6615_ ( .A(\RegFile/_2524_ ), .B1(\RegFile/_3519_ ), .B2(\RegFile/_2047_ ), .C1(\RegFile/_3295_ ), .C2(\RegFile/_2121_ ), .ZN(\RegFile/_2525_ ) );
NAND3_X1 \RegFile/_6616_ ( .A1(\RegFile/_2012_ ), .A2(\RegFile/_3423_ ), .A3(\RegFile/_1994_ ), .ZN(\RegFile/_2526_ ) );
NAND3_X1 \RegFile/_6617_ ( .A1(\RegFile/_1994_ ), .A2(\RegFile/_2003_ ), .A3(\RegFile/_3391_ ), .ZN(\RegFile/_2527_ ) );
NAND2_X1 \RegFile/_6618_ ( .A1(\RegFile/_2526_ ), .A2(\RegFile/_2527_ ), .ZN(\RegFile/_2528_ ) );
AOI221_X4 \RegFile/_6619_ ( .A(\RegFile/_2528_ ), .B1(\RegFile/_3359_ ), .B2(\RegFile/_2126_ ), .C1(\RegFile/_3327_ ), .C2(\RegFile/_2127_ ), .ZN(\RegFile/_2529_ ) );
NAND4_X4 \RegFile/_6620_ ( .A1(\RegFile/_2522_ ), .A2(\RegFile/_2062_ ), .A3(\RegFile/_2525_ ), .A4(\RegFile/_2529_ ), .ZN(\RegFile/_2530_ ) );
OR3_X1 \RegFile/_6621_ ( .A1(\RegFile/_2066_ ), .A2(\RegFile/_2068_ ), .A3(\RegFile/_0729_ ), .ZN(\RegFile/_2531_ ) );
NAND2_X1 \RegFile/_6622_ ( .A1(\RegFile/_2530_ ), .A2(\RegFile/_2531_ ), .ZN(\RegFile/_2532_ ) );
BUF_X4 \RegFile/_6623_ ( .A(\RegFile/_2532_ ), .Z(\RegFile/_2533_ ) );
AOI21_X1 \RegFile/_6624_ ( .A(\RegFile/_2515_ ), .B1(\RegFile/_2533_ ), .B2(\RegFile/_2400_ ), .ZN(\RegFile/_0629_ ) );
NAND2_X1 \RegFile/_6625_ ( .A1(\RegFile/_2077_ ), .A2(\RegFile/_3488_ ), .ZN(\RegFile/_2534_ ) );
NAND3_X1 \RegFile/_6626_ ( .A1(\RegFile/_2090_ ), .A2(\RegFile/_3552_ ), .A3(\RegFile/_2091_ ), .ZN(\RegFile/_2535_ ) );
OAI21_X1 \RegFile/_6627_ ( .A(\RegFile/_2535_ ), .B1(\RegFile/_2145_ ), .B2(\RegFile/_1833_ ), .ZN(\RegFile/_2536_ ) );
AOI221_X4 \RegFile/_6628_ ( .A(\RegFile/_2536_ ), .B1(\RegFile/_3648_ ), .B2(\RegFile/_2044_ ), .C1(\RegFile/_3616_ ), .C2(\RegFile/_2053_ ), .ZN(\RegFile/_2537_ ) );
AOI22_X1 \RegFile/_6629_ ( .A1(\RegFile/_2048_ ), .A2(\RegFile/_3520_ ), .B1(\RegFile/_3296_ ), .B2(\RegFile/_2083_ ), .ZN(\RegFile/_2538_ ) );
AOI22_X1 \RegFile/_6630_ ( .A1(\RegFile/_3328_ ), .A2(\RegFile/_2127_ ), .B1(\RegFile/_2081_ ), .B2(\RegFile/_3360_ ), .ZN(\RegFile/_2539_ ) );
AND3_X1 \RegFile/_6631_ ( .A1(\RegFile/_2220_ ), .A2(\RegFile/_2090_ ), .A3(\RegFile/_3680_ ), .ZN(\RegFile/_2540_ ) );
AOI21_X1 \RegFile/_6632_ ( .A(\RegFile/_2540_ ), .B1(\RegFile/_3712_ ), .B2(\RegFile/_2009_ ), .ZN(\RegFile/_2541_ ) );
AOI22_X1 \RegFile/_6633_ ( .A1(\RegFile/_2085_ ), .A2(\RegFile/_3424_ ), .B1(\RegFile/_3392_ ), .B2(\RegFile/_2086_ ), .ZN(\RegFile/_2542_ ) );
AND4_X1 \RegFile/_6634_ ( .A1(\RegFile/_2538_ ), .A2(\RegFile/_2539_ ), .A3(\RegFile/_2541_ ), .A4(\RegFile/_2542_ ), .ZN(\RegFile/_2543_ ) );
NAND3_X1 \RegFile/_6635_ ( .A1(\RegFile/_2096_ ), .A2(\RegFile/_2098_ ), .A3(\RegFile/_3776_ ), .ZN(\RegFile/_2544_ ) );
NAND3_X1 \RegFile/_6636_ ( .A1(\RegFile/_2268_ ), .A2(\RegFile/_3744_ ), .A3(\RegFile/_2101_ ), .ZN(\RegFile/_2545_ ) );
NAND3_X1 \RegFile/_6637_ ( .A1(\RegFile/_1989_ ), .A2(\RegFile/_2255_ ), .A3(\RegFile/_3488_ ), .ZN(\RegFile/_2546_ ) );
NAND3_X1 \RegFile/_6638_ ( .A1(\RegFile/_2107_ ), .A2(\RegFile/_3456_ ), .A3(\RegFile/_2104_ ), .ZN(\RegFile/_2547_ ) );
AND4_X1 \RegFile/_6639_ ( .A1(\RegFile/_2544_ ), .A2(\RegFile/_2545_ ), .A3(\RegFile/_2546_ ), .A4(\RegFile/_2547_ ), .ZN(\RegFile/_2548_ ) );
NAND4_X1 \RegFile/_6640_ ( .A1(\RegFile/_2537_ ), .A2(\RegFile/_2089_ ), .A3(\RegFile/_2543_ ), .A4(\RegFile/_2548_ ), .ZN(\RegFile/_2549_ ) );
OR3_X1 \RegFile/_6641_ ( .A1(\RegFile/_2236_ ), .A2(\RegFile/_2237_ ), .A3(\RegFile/_0730_ ), .ZN(\RegFile/_2550_ ) );
NAND2_X1 \RegFile/_6642_ ( .A1(\RegFile/_2549_ ), .A2(\RegFile/_2550_ ), .ZN(\RegFile/_2551_ ) );
BUF_X4 \RegFile/_6643_ ( .A(\RegFile/_2551_ ), .Z(\RegFile/_2552_ ) );
OAI21_X1 \RegFile/_6644_ ( .A(\RegFile/_2534_ ), .B1(\RegFile/_2552_ ), .B2(\RegFile/_2114_ ), .ZN(\RegFile/_0630_ ) );
AOI21_X1 \RegFile/_6645_ ( .A(\RegFile/_3489_ ), .B1(\RegFile/_2380_ ), .B2(\RegFile/_2357_ ), .ZN(\RegFile/_2553_ ) );
NAND3_X1 \RegFile/_6646_ ( .A1(\RegFile/_2090_ ), .A2(\RegFile/_3553_ ), .A3(\RegFile/_2091_ ), .ZN(\RegFile/_2554_ ) );
OAI21_X1 \RegFile/_6647_ ( .A(\RegFile/_2554_ ), .B1(\RegFile/_2145_ ), .B2(\RegFile/_1853_ ), .ZN(\RegFile/_2555_ ) );
AOI221_X4 \RegFile/_6648_ ( .A(\RegFile/_2555_ ), .B1(\RegFile/_3649_ ), .B2(\RegFile/_2044_ ), .C1(\RegFile/_3617_ ), .C2(\RegFile/_2053_ ), .ZN(\RegFile/_2556_ ) );
AOI22_X1 \RegFile/_6649_ ( .A1(\RegFile/_2048_ ), .A2(\RegFile/_3521_ ), .B1(\RegFile/_3297_ ), .B2(\RegFile/_2083_ ), .ZN(\RegFile/_2557_ ) );
AOI22_X1 \RegFile/_6650_ ( .A1(\RegFile/_3329_ ), .A2(\RegFile/_2127_ ), .B1(\RegFile/_2081_ ), .B2(\RegFile/_3361_ ), .ZN(\RegFile/_2558_ ) );
AND3_X1 \RegFile/_6651_ ( .A1(\RegFile/_2220_ ), .A2(\RegFile/_2090_ ), .A3(\RegFile/_3681_ ), .ZN(\RegFile/_2559_ ) );
AOI21_X1 \RegFile/_6652_ ( .A(\RegFile/_2559_ ), .B1(\RegFile/_3713_ ), .B2(\RegFile/_2009_ ), .ZN(\RegFile/_2560_ ) );
AOI22_X1 \RegFile/_6653_ ( .A1(\RegFile/_2085_ ), .A2(\RegFile/_3425_ ), .B1(\RegFile/_3393_ ), .B2(\RegFile/_2086_ ), .ZN(\RegFile/_2561_ ) );
AND4_X1 \RegFile/_6654_ ( .A1(\RegFile/_2557_ ), .A2(\RegFile/_2558_ ), .A3(\RegFile/_2560_ ), .A4(\RegFile/_2561_ ), .ZN(\RegFile/_2562_ ) );
NAND3_X1 \RegFile/_6655_ ( .A1(\RegFile/_2096_ ), .A2(\RegFile/_2098_ ), .A3(\RegFile/_3777_ ), .ZN(\RegFile/_2563_ ) );
NAND3_X1 \RegFile/_6656_ ( .A1(\RegFile/_2268_ ), .A2(\RegFile/_3745_ ), .A3(\RegFile/_2101_ ), .ZN(\RegFile/_2564_ ) );
NAND3_X1 \RegFile/_6657_ ( .A1(\RegFile/_1989_ ), .A2(\RegFile/_2255_ ), .A3(\RegFile/_3489_ ), .ZN(\RegFile/_2565_ ) );
NAND3_X1 \RegFile/_6658_ ( .A1(\RegFile/_2107_ ), .A2(\RegFile/_3457_ ), .A3(\RegFile/_2104_ ), .ZN(\RegFile/_2566_ ) );
AND4_X1 \RegFile/_6659_ ( .A1(\RegFile/_2563_ ), .A2(\RegFile/_2564_ ), .A3(\RegFile/_2565_ ), .A4(\RegFile/_2566_ ), .ZN(\RegFile/_2567_ ) );
NAND4_X1 \RegFile/_6660_ ( .A1(\RegFile/_2556_ ), .A2(\RegFile/_2089_ ), .A3(\RegFile/_2562_ ), .A4(\RegFile/_2567_ ), .ZN(\RegFile/_2568_ ) );
OR3_X1 \RegFile/_6661_ ( .A1(\RegFile/_2236_ ), .A2(\RegFile/_2237_ ), .A3(\RegFile/_0731_ ), .ZN(\RegFile/_2569_ ) );
NAND2_X1 \RegFile/_6662_ ( .A1(\RegFile/_2568_ ), .A2(\RegFile/_2569_ ), .ZN(\RegFile/_2570_ ) );
BUF_X4 \RegFile/_6663_ ( .A(\RegFile/_2570_ ), .Z(\RegFile/_2571_ ) );
AOI21_X1 \RegFile/_6664_ ( .A(\RegFile/_2553_ ), .B1(\RegFile/_2571_ ), .B2(\RegFile/_2400_ ), .ZN(\RegFile/_0631_ ) );
NAND2_X1 \RegFile/_6665_ ( .A1(\RegFile/_2077_ ), .A2(\RegFile/_3490_ ), .ZN(\RegFile/_2572_ ) );
NAND3_X1 \RegFile/_6666_ ( .A1(\RegFile/_2161_ ), .A2(\RegFile/_3650_ ), .A3(\RegFile/_2338_ ), .ZN(\RegFile/_2573_ ) );
AND3_X1 \RegFile/_6667_ ( .A1(\RegFile/_2026_ ), .A2(\RegFile/_3554_ ), .A3(\RegFile/_2037_ ), .ZN(\RegFile/_2574_ ) );
AOI221_X1 \RegFile/_6668_ ( .A(\RegFile/_2574_ ), .B1(\RegFile/_3298_ ), .B2(\RegFile/_2059_ ), .C1(\RegFile/_3522_ ), .C2(\RegFile/_2047_ ), .ZN(\RegFile/_2575_ ) );
NAND3_X1 \RegFile/_6669_ ( .A1(\RegFile/_2338_ ), .A2(\RegFile/_2254_ ), .A3(\RegFile/_3682_ ), .ZN(\RegFile/_2576_ ) );
AOI22_X1 \RegFile/_6670_ ( .A1(\RegFile/_2053_ ), .A2(\RegFile/_3618_ ), .B1(\RegFile/_2055_ ), .B2(\RegFile/_3586_ ), .ZN(\RegFile/_2577_ ) );
AND4_X1 \RegFile/_6671_ ( .A1(\RegFile/_2573_ ), .A2(\RegFile/_2575_ ), .A3(\RegFile/_2576_ ), .A4(\RegFile/_2577_ ), .ZN(\RegFile/_2578_ ) );
NAND3_X1 \RegFile/_6672_ ( .A1(\RegFile/_1990_ ), .A2(\RegFile/_1996_ ), .A3(\RegFile/_3490_ ), .ZN(\RegFile/_2579_ ) );
NAND3_X1 \RegFile/_6673_ ( .A1(\RegFile/_2096_ ), .A2(\RegFile/_2098_ ), .A3(\RegFile/_3778_ ), .ZN(\RegFile/_2580_ ) );
NAND3_X1 \RegFile/_6674_ ( .A1(\RegFile/_2097_ ), .A2(\RegFile/_3426_ ), .A3(\RegFile/_2103_ ), .ZN(\RegFile/_2581_ ) );
NAND3_X1 \RegFile/_6675_ ( .A1(\RegFile/_2001_ ), .A2(\RegFile/_3362_ ), .A3(\RegFile/_1988_ ), .ZN(\RegFile/_2582_ ) );
NAND3_X1 \RegFile/_6676_ ( .A1(\RegFile/_2041_ ), .A2(\RegFile/_3458_ ), .A3(\RegFile/_2103_ ), .ZN(\RegFile/_2583_ ) );
NAND3_X1 \RegFile/_6677_ ( .A1(\RegFile/_2103_ ), .A2(\RegFile/_2034_ ), .A3(\RegFile/_3394_ ), .ZN(\RegFile/_2584_ ) );
AND4_X1 \RegFile/_6678_ ( .A1(\RegFile/_2581_ ), .A2(\RegFile/_2582_ ), .A3(\RegFile/_2583_ ), .A4(\RegFile/_2584_ ), .ZN(\RegFile/_2585_ ) );
NAND3_X1 \RegFile/_6679_ ( .A1(\RegFile/_2100_ ), .A2(\RegFile/_3330_ ), .A3(\RegFile/_2107_ ), .ZN(\RegFile/_2586_ ) );
AOI22_X1 \RegFile/_6680_ ( .A1(\RegFile/_2131_ ), .A2(\RegFile/_3746_ ), .B1(\RegFile/_2008_ ), .B2(\RegFile/_3714_ ), .ZN(\RegFile/_2587_ ) );
AND4_X1 \RegFile/_6681_ ( .A1(\RegFile/_2580_ ), .A2(\RegFile/_2585_ ), .A3(\RegFile/_2586_ ), .A4(\RegFile/_2587_ ), .ZN(\RegFile/_2588_ ) );
NAND4_X1 \RegFile/_6682_ ( .A1(\RegFile/_2578_ ), .A2(\RegFile/_2089_ ), .A3(\RegFile/_2579_ ), .A4(\RegFile/_2588_ ), .ZN(\RegFile/_2589_ ) );
OR3_X1 \RegFile/_6683_ ( .A1(\RegFile/_2236_ ), .A2(\RegFile/_2237_ ), .A3(\RegFile/_0732_ ), .ZN(\RegFile/_2590_ ) );
NAND2_X1 \RegFile/_6684_ ( .A1(\RegFile/_2589_ ), .A2(\RegFile/_2590_ ), .ZN(\RegFile/_2591_ ) );
BUF_X4 \RegFile/_6685_ ( .A(\RegFile/_2591_ ), .Z(\RegFile/_2592_ ) );
OAI21_X1 \RegFile/_6686_ ( .A(\RegFile/_2572_ ), .B1(\RegFile/_2592_ ), .B2(\RegFile/_2114_ ), .ZN(\RegFile/_0632_ ) );
NAND2_X1 \RegFile/_6687_ ( .A1(\RegFile/_2077_ ), .A2(\RegFile/_3491_ ), .ZN(\RegFile/_2593_ ) );
OAI22_X1 \RegFile/_6688_ ( .A1(\RegFile/_2144_ ), .A2(\RegFile/_1272_ ), .B1(\RegFile/_2146_ ), .B2(\RegFile/_1271_ ), .ZN(\RegFile/_2594_ ) );
AOI221_X4 \RegFile/_6689_ ( .A(\RegFile/_2594_ ), .B1(\RegFile/_3651_ ), .B2(\RegFile/_2133_ ), .C1(\RegFile/_3619_ ), .C2(\RegFile/_2149_ ), .ZN(\RegFile/_2595_ ) );
AND3_X1 \RegFile/_6690_ ( .A1(\RegFile/_2040_ ), .A2(\RegFile/_2168_ ), .A3(\RegFile/_3683_ ), .ZN(\RegFile/_2596_ ) );
AOI21_X1 \RegFile/_6691_ ( .A(\RegFile/_2596_ ), .B1(\RegFile/_3715_ ), .B2(\RegFile/_2152_ ), .ZN(\RegFile/_2597_ ) );
AOI22_X1 \RegFile/_6692_ ( .A1(\RegFile/_3331_ ), .A2(\RegFile/_2018_ ), .B1(\RegFile/_2021_ ), .B2(\RegFile/_3363_ ), .ZN(\RegFile/_2598_ ) );
AOI22_X1 \RegFile/_6693_ ( .A1(\RegFile/_2155_ ), .A2(\RegFile/_3523_ ), .B1(\RegFile/_3299_ ), .B2(\RegFile/_2121_ ), .ZN(\RegFile/_2599_ ) );
AOI22_X1 \RegFile/_6694_ ( .A1(\RegFile/_2031_ ), .A2(\RegFile/_3427_ ), .B1(\RegFile/_3395_ ), .B2(\RegFile/_2024_ ), .ZN(\RegFile/_2600_ ) );
AND4_X1 \RegFile/_6695_ ( .A1(\RegFile/_2597_ ), .A2(\RegFile/_2598_ ), .A3(\RegFile/_2599_ ), .A4(\RegFile/_2600_ ), .ZN(\RegFile/_2601_ ) );
NAND3_X1 \RegFile/_6696_ ( .A1(\RegFile/_2027_ ), .A2(\RegFile/_3459_ ), .A3(\RegFile/_2028_ ), .ZN(\RegFile/_2602_ ) );
NAND3_X1 \RegFile/_6697_ ( .A1(\RegFile/_2165_ ), .A2(\RegFile/_2028_ ), .A3(\RegFile/_3491_ ), .ZN(\RegFile/_2603_ ) );
NAND2_X1 \RegFile/_6698_ ( .A1(\RegFile/_2602_ ), .A2(\RegFile/_2603_ ), .ZN(\RegFile/_2604_ ) );
AOI221_X4 \RegFile/_6699_ ( .A(\RegFile/_2604_ ), .B1(\RegFile/_2130_ ), .B2(\RegFile/_3779_ ), .C1(\RegFile/_3747_ ), .C2(\RegFile/_2131_ ), .ZN(\RegFile/_2605_ ) );
NAND4_X4 \RegFile/_6700_ ( .A1(\RegFile/_2595_ ), .A2(\RegFile/_2063_ ), .A3(\RegFile/_2601_ ), .A4(\RegFile/_2605_ ), .ZN(\RegFile/_2606_ ) );
OR3_X2 \RegFile/_6701_ ( .A1(\RegFile/_2067_ ), .A2(\RegFile/_2069_ ), .A3(\RegFile/_0733_ ), .ZN(\RegFile/_2607_ ) );
NAND2_X2 \RegFile/_6702_ ( .A1(\RegFile/_2606_ ), .A2(\RegFile/_2607_ ), .ZN(\RegFile/_2608_ ) );
OAI21_X1 \RegFile/_6703_ ( .A(\RegFile/_2593_ ), .B1(\RegFile/_2608_ ), .B2(\RegFile/_2114_ ), .ZN(\RegFile/_0633_ ) );
AOI21_X1 \RegFile/_6704_ ( .A(\RegFile/_3492_ ), .B1(\RegFile/_2380_ ), .B2(\RegFile/_2357_ ), .ZN(\RegFile/_2609_ ) );
AND3_X1 \RegFile/_6705_ ( .A1(\RegFile/_2040_ ), .A2(\RegFile/_2027_ ), .A3(\RegFile/_3684_ ), .ZN(\RegFile/_2610_ ) );
AOI21_X1 \RegFile/_6706_ ( .A(\RegFile/_2610_ ), .B1(\RegFile/_3716_ ), .B2(\RegFile/_2152_ ), .ZN(\RegFile/_2611_ ) );
AOI22_X1 \RegFile/_6707_ ( .A1(\RegFile/_3332_ ), .A2(\RegFile/_2018_ ), .B1(\RegFile/_2081_ ), .B2(\RegFile/_3364_ ), .ZN(\RegFile/_2612_ ) );
AOI22_X1 \RegFile/_6708_ ( .A1(\RegFile/_2048_ ), .A2(\RegFile/_3524_ ), .B1(\RegFile/_3300_ ), .B2(\RegFile/_2121_ ), .ZN(\RegFile/_2613_ ) );
AOI22_X1 \RegFile/_6709_ ( .A1(\RegFile/_2085_ ), .A2(\RegFile/_3428_ ), .B1(\RegFile/_3396_ ), .B2(\RegFile/_2086_ ), .ZN(\RegFile/_2614_ ) );
AND4_X1 \RegFile/_6710_ ( .A1(\RegFile/_2611_ ), .A2(\RegFile/_2612_ ), .A3(\RegFile/_2613_ ), .A4(\RegFile/_2614_ ), .ZN(\RegFile/_2615_ ) );
NAND3_X1 \RegFile/_6711_ ( .A1(\RegFile/_2041_ ), .A2(\RegFile/_3556_ ), .A3(\RegFile/_2091_ ), .ZN(\RegFile/_2616_ ) );
NAND3_X1 \RegFile/_6712_ ( .A1(\RegFile/_1988_ ), .A2(\RegFile/_2091_ ), .A3(\RegFile/_3588_ ), .ZN(\RegFile/_2617_ ) );
NAND2_X1 \RegFile/_6713_ ( .A1(\RegFile/_2616_ ), .A2(\RegFile/_2617_ ), .ZN(\RegFile/_2618_ ) );
AOI221_X4 \RegFile/_6714_ ( .A(\RegFile/_2618_ ), .B1(\RegFile/_3620_ ), .B2(\RegFile/_2134_ ), .C1(\RegFile/_3652_ ), .C2(\RegFile/_2133_ ), .ZN(\RegFile/_2619_ ) );
NAND3_X1 \RegFile/_6715_ ( .A1(\RegFile/_2096_ ), .A2(\RegFile/_2161_ ), .A3(\RegFile/_3780_ ), .ZN(\RegFile/_2620_ ) );
NAND3_X1 \RegFile/_6716_ ( .A1(\RegFile/_2268_ ), .A2(\RegFile/_3748_ ), .A3(\RegFile/_2163_ ), .ZN(\RegFile/_2621_ ) );
NAND3_X1 \RegFile/_6717_ ( .A1(\RegFile/_2166_ ), .A2(\RegFile/_2255_ ), .A3(\RegFile/_3492_ ), .ZN(\RegFile/_2622_ ) );
NAND3_X1 \RegFile/_6718_ ( .A1(\RegFile/_2254_ ), .A2(\RegFile/_3460_ ), .A3(\RegFile/_2255_ ), .ZN(\RegFile/_2623_ ) );
AND4_X1 \RegFile/_6719_ ( .A1(\RegFile/_2620_ ), .A2(\RegFile/_2621_ ), .A3(\RegFile/_2622_ ), .A4(\RegFile/_2623_ ), .ZN(\RegFile/_2624_ ) );
NAND4_X1 \RegFile/_6720_ ( .A1(\RegFile/_2615_ ), .A2(\RegFile/_2063_ ), .A3(\RegFile/_2619_ ), .A4(\RegFile/_2624_ ), .ZN(\RegFile/_2625_ ) );
OR3_X1 \RegFile/_6721_ ( .A1(\RegFile/_2236_ ), .A2(\RegFile/_2237_ ), .A3(\RegFile/_0734_ ), .ZN(\RegFile/_2626_ ) );
NAND2_X1 \RegFile/_6722_ ( .A1(\RegFile/_2625_ ), .A2(\RegFile/_2626_ ), .ZN(\RegFile/_2627_ ) );
BUF_X4 \RegFile/_6723_ ( .A(\RegFile/_2627_ ), .Z(\RegFile/_2628_ ) );
AOI21_X1 \RegFile/_6724_ ( .A(\RegFile/_2609_ ), .B1(\RegFile/_2628_ ), .B2(\RegFile/_2400_ ), .ZN(\RegFile/_0634_ ) );
AOI21_X1 \RegFile/_6725_ ( .A(\RegFile/_3493_ ), .B1(\RegFile/_2380_ ), .B2(\RegFile/_2357_ ), .ZN(\RegFile/_2629_ ) );
NAND3_X1 \RegFile/_6726_ ( .A1(\RegFile/_2090_ ), .A2(\RegFile/_3557_ ), .A3(\RegFile/_2037_ ), .ZN(\RegFile/_2630_ ) );
OAI21_X1 \RegFile/_6727_ ( .A(\RegFile/_2630_ ), .B1(\RegFile/_2145_ ), .B2(\RegFile/_1912_ ), .ZN(\RegFile/_2631_ ) );
AOI221_X4 \RegFile/_6728_ ( .A(\RegFile/_2631_ ), .B1(\RegFile/_3653_ ), .B2(\RegFile/_2044_ ), .C1(\RegFile/_3621_ ), .C2(\RegFile/_2053_ ), .ZN(\RegFile/_2632_ ) );
AOI22_X1 \RegFile/_6729_ ( .A1(\RegFile/_2048_ ), .A2(\RegFile/_3525_ ), .B1(\RegFile/_3301_ ), .B2(\RegFile/_2083_ ), .ZN(\RegFile/_2633_ ) );
AOI22_X1 \RegFile/_6730_ ( .A1(\RegFile/_3333_ ), .A2(\RegFile/_2127_ ), .B1(\RegFile/_2126_ ), .B2(\RegFile/_3365_ ), .ZN(\RegFile/_2634_ ) );
AND3_X1 \RegFile/_6731_ ( .A1(\RegFile/_2220_ ), .A2(\RegFile/_2106_ ), .A3(\RegFile/_3685_ ), .ZN(\RegFile/_2635_ ) );
AOI21_X1 \RegFile/_6732_ ( .A(\RegFile/_2635_ ), .B1(\RegFile/_3717_ ), .B2(\RegFile/_2009_ ), .ZN(\RegFile/_2636_ ) );
AOI22_X1 \RegFile/_6733_ ( .A1(\RegFile/_2188_ ), .A2(\RegFile/_3429_ ), .B1(\RegFile/_3397_ ), .B2(\RegFile/_2023_ ), .ZN(\RegFile/_2637_ ) );
AND4_X1 \RegFile/_6734_ ( .A1(\RegFile/_2633_ ), .A2(\RegFile/_2634_ ), .A3(\RegFile/_2636_ ), .A4(\RegFile/_2637_ ), .ZN(\RegFile/_2638_ ) );
AOI22_X1 \RegFile/_6735_ ( .A1(\RegFile/_3781_ ), .A2(\RegFile/_2014_ ), .B1(\RegFile/_2131_ ), .B2(\RegFile/_3749_ ), .ZN(\RegFile/_2639_ ) );
NAND3_X1 \RegFile/_6736_ ( .A1(\RegFile/_2166_ ), .A2(\RegFile/_2170_ ), .A3(\RegFile/_3493_ ), .ZN(\RegFile/_2640_ ) );
NAND3_X1 \RegFile/_6737_ ( .A1(\RegFile/_2254_ ), .A2(\RegFile/_3461_ ), .A3(\RegFile/_2170_ ), .ZN(\RegFile/_2641_ ) );
AND3_X1 \RegFile/_6738_ ( .A1(\RegFile/_2639_ ), .A2(\RegFile/_2640_ ), .A3(\RegFile/_2641_ ), .ZN(\RegFile/_2642_ ) );
NAND4_X1 \RegFile/_6739_ ( .A1(\RegFile/_2632_ ), .A2(\RegFile/_2089_ ), .A3(\RegFile/_2638_ ), .A4(\RegFile/_2642_ ), .ZN(\RegFile/_2643_ ) );
OR3_X1 \RegFile/_6740_ ( .A1(\RegFile/_2066_ ), .A2(\RegFile/_2068_ ), .A3(\RegFile/_0735_ ), .ZN(\RegFile/_2644_ ) );
NAND2_X1 \RegFile/_6741_ ( .A1(\RegFile/_2643_ ), .A2(\RegFile/_2644_ ), .ZN(\RegFile/_2645_ ) );
BUF_X4 \RegFile/_6742_ ( .A(\RegFile/_2645_ ), .Z(\RegFile/_2646_ ) );
AOI21_X1 \RegFile/_6743_ ( .A(\RegFile/_2629_ ), .B1(\RegFile/_2646_ ), .B2(\RegFile/_2400_ ), .ZN(\RegFile/_0635_ ) );
NAND2_X1 \RegFile/_6744_ ( .A1(\RegFile/_2076_ ), .A2(\RegFile/_3494_ ), .ZN(\RegFile/_2647_ ) );
NAND3_X1 \RegFile/_6745_ ( .A1(\RegFile/_2006_ ), .A2(\RegFile/_3622_ ), .A3(\RegFile/_2003_ ), .ZN(\RegFile/_2648_ ) );
OAI21_X2 \RegFile/_6746_ ( .A(\RegFile/_2648_ ), .B1(\RegFile/_2181_ ), .B2(\RegFile/_1315_ ), .ZN(\RegFile/_2649_ ) );
AOI221_X2 \RegFile/_6747_ ( .A(\RegFile/_2649_ ), .B1(\RegFile/_3590_ ), .B2(\RegFile/_2054_ ), .C1(\RegFile/_3558_ ), .C2(\RegFile/_2049_ ), .ZN(\RegFile/_2650_ ) );
NAND3_X1 \RegFile/_6748_ ( .A1(\RegFile/_1989_ ), .A2(\RegFile/_2104_ ), .A3(\RegFile/_3494_ ), .ZN(\RegFile/_2651_ ) );
NAND3_X1 \RegFile/_6749_ ( .A1(\RegFile/_2107_ ), .A2(\RegFile/_3462_ ), .A3(\RegFile/_2104_ ), .ZN(\RegFile/_2652_ ) );
AOI22_X1 \RegFile/_6750_ ( .A1(\RegFile/_3782_ ), .A2(\RegFile/_2130_ ), .B1(\RegFile/_2004_ ), .B2(\RegFile/_3750_ ), .ZN(\RegFile/_2653_ ) );
NAND4_X1 \RegFile/_6751_ ( .A1(\RegFile/_2650_ ), .A2(\RegFile/_2651_ ), .A3(\RegFile/_2652_ ), .A4(\RegFile/_2653_ ), .ZN(\RegFile/_2654_ ) );
AOI22_X1 \RegFile/_6752_ ( .A1(\RegFile/_2047_ ), .A2(\RegFile/_3526_ ), .B1(\RegFile/_3302_ ), .B2(\RegFile/_2059_ ), .ZN(\RegFile/_2655_ ) );
OAI221_X1 \RegFile/_6753_ ( .A(\RegFile/_2655_ ), .B1(\RegFile/_1318_ ), .B2(\RegFile/_2116_ ), .C1(\RegFile/_1314_ ), .C2(\RegFile/_2118_ ), .ZN(\RegFile/_2656_ ) );
AOI22_X1 \RegFile/_6754_ ( .A1(\RegFile/_2188_ ), .A2(\RegFile/_3430_ ), .B1(\RegFile/_3398_ ), .B2(\RegFile/_2023_ ), .ZN(\RegFile/_2657_ ) );
NAND3_X1 \RegFile/_6755_ ( .A1(\RegFile/_2159_ ), .A2(\RegFile/_3334_ ), .A3(\RegFile/_2168_ ), .ZN(\RegFile/_2658_ ) );
NAND3_X1 \RegFile/_6756_ ( .A1(\RegFile/_2159_ ), .A2(\RegFile/_3366_ ), .A3(\RegFile/_2165_ ), .ZN(\RegFile/_2659_ ) );
NAND3_X1 \RegFile/_6757_ ( .A1(\RegFile/_2657_ ), .A2(\RegFile/_2658_ ), .A3(\RegFile/_2659_ ), .ZN(\RegFile/_2660_ ) );
NOR4_X2 \RegFile/_6758_ ( .A1(\RegFile/_2654_ ), .A2(\RegFile/_2061_ ), .A3(\RegFile/_2656_ ), .A4(\RegFile/_2660_ ), .ZN(\RegFile/_2661_ ) );
AOI211_X4 \RegFile/_6759_ ( .A(\RegFile/_2060_ ), .B(\RegFile/_0736_ ), .C1(\RegFile/_2163_ ), .C2(\RegFile/_2038_ ), .ZN(\RegFile/_2662_ ) );
OR2_X4 \RegFile/_6760_ ( .A1(\RegFile/_2661_ ), .A2(\RegFile/_2662_ ), .ZN(\RegFile/_2663_ ) );
BUF_X8 \RegFile/_6761_ ( .A(\RegFile/_2663_ ), .Z(\RegFile/_2664_ ) );
OAI21_X1 \RegFile/_6762_ ( .A(\RegFile/_2647_ ), .B1(\RegFile/_2664_ ), .B2(\RegFile/_2114_ ), .ZN(\RegFile/_0636_ ) );
BUF_X4 \RegFile/_6763_ ( .A(\RegFile/_1996_ ), .Z(\RegFile/_2665_ ) );
AOI21_X1 \RegFile/_6764_ ( .A(\RegFile/_3495_ ), .B1(\RegFile/_2380_ ), .B2(\RegFile/_2665_ ), .ZN(\RegFile/_2666_ ) );
AOI22_X1 \RegFile/_6765_ ( .A1(\RegFile/_2045_ ), .A2(\RegFile/_3655_ ), .B1(\RegFile/_2134_ ), .B2(\RegFile/_3623_ ), .ZN(\RegFile/_2667_ ) );
INV_X1 \RegFile/_6766_ ( .A(\RegFile/_3591_ ), .ZN(\RegFile/_2668_ ) );
INV_X1 \RegFile/_6767_ ( .A(\RegFile/_3559_ ), .ZN(\RegFile/_2669_ ) );
OAI221_X1 \RegFile/_6768_ ( .A(\RegFile/_2667_ ), .B1(\RegFile/_2668_ ), .B2(\RegFile/_2146_ ), .C1(\RegFile/_2669_ ), .C2(\RegFile/_2144_ ), .ZN(\RegFile/_2670_ ) );
AOI22_X1 \RegFile/_6769_ ( .A1(\RegFile/_3335_ ), .A2(\RegFile/_2127_ ), .B1(\RegFile/_2126_ ), .B2(\RegFile/_3367_ ), .ZN(\RegFile/_2671_ ) );
AND3_X1 \RegFile/_6770_ ( .A1(\RegFile/_2117_ ), .A2(\RegFile/_2106_ ), .A3(\RegFile/_3687_ ), .ZN(\RegFile/_2672_ ) );
AOI21_X1 \RegFile/_6771_ ( .A(\RegFile/_2672_ ), .B1(\RegFile/_3719_ ), .B2(\RegFile/_2008_ ), .ZN(\RegFile/_2673_ ) );
AOI22_X1 \RegFile/_6772_ ( .A1(\RegFile/_2120_ ), .A2(\RegFile/_3527_ ), .B1(\RegFile/_3303_ ), .B2(\RegFile/_2083_ ), .ZN(\RegFile/_2674_ ) );
AOI22_X1 \RegFile/_6773_ ( .A1(\RegFile/_2188_ ), .A2(\RegFile/_3431_ ), .B1(\RegFile/_3399_ ), .B2(\RegFile/_2023_ ), .ZN(\RegFile/_2675_ ) );
NAND4_X1 \RegFile/_6774_ ( .A1(\RegFile/_2671_ ), .A2(\RegFile/_2673_ ), .A3(\RegFile/_2674_ ), .A4(\RegFile/_2675_ ), .ZN(\RegFile/_2676_ ) );
NAND3_X1 \RegFile/_6775_ ( .A1(\RegFile/_2100_ ), .A2(\RegFile/_2098_ ), .A3(\RegFile/_3783_ ), .ZN(\RegFile/_2677_ ) );
NAND3_X1 \RegFile/_6776_ ( .A1(\RegFile/_2100_ ), .A2(\RegFile/_3751_ ), .A3(\RegFile/_2101_ ), .ZN(\RegFile/_2678_ ) );
NAND3_X1 \RegFile/_6777_ ( .A1(\RegFile/_1989_ ), .A2(\RegFile/_2104_ ), .A3(\RegFile/_3495_ ), .ZN(\RegFile/_2679_ ) );
NAND3_X1 \RegFile/_6778_ ( .A1(\RegFile/_2107_ ), .A2(\RegFile/_3463_ ), .A3(\RegFile/_1995_ ), .ZN(\RegFile/_2680_ ) );
NAND4_X1 \RegFile/_6779_ ( .A1(\RegFile/_2677_ ), .A2(\RegFile/_2678_ ), .A3(\RegFile/_2679_ ), .A4(\RegFile/_2680_ ), .ZN(\RegFile/_2681_ ) );
NOR4_X2 \RegFile/_6780_ ( .A1(\RegFile/_2670_ ), .A2(\RegFile/_2676_ ), .A3(\RegFile/_2061_ ), .A4(\RegFile/_2681_ ), .ZN(\RegFile/_2682_ ) );
AOI211_X4 \RegFile/_6781_ ( .A(\RegFile/_2068_ ), .B(\RegFile/_0737_ ), .C1(\RegFile/_2035_ ), .C2(\RegFile/_2376_ ), .ZN(\RegFile/_2683_ ) );
OR2_X2 \RegFile/_6782_ ( .A1(\RegFile/_2682_ ), .A2(\RegFile/_2683_ ), .ZN(\RegFile/_2684_ ) );
BUF_X4 \RegFile/_6783_ ( .A(\RegFile/_2684_ ), .Z(\RegFile/_2685_ ) );
AOI21_X1 \RegFile/_6784_ ( .A(\RegFile/_2666_ ), .B1(\RegFile/_2685_ ), .B2(\RegFile/_2400_ ), .ZN(\RegFile/_0637_ ) );
NAND2_X1 \RegFile/_6785_ ( .A1(\RegFile/_2076_ ), .A2(\RegFile/_3497_ ), .ZN(\RegFile/_2686_ ) );
NAND3_X1 \RegFile/_6786_ ( .A1(\RegFile/_2041_ ), .A2(\RegFile/_3561_ ), .A3(\RegFile/_2091_ ), .ZN(\RegFile/_2687_ ) );
INV_X1 \RegFile/_6787_ ( .A(\RegFile/_3593_ ), .ZN(\RegFile/_2688_ ) );
OAI21_X1 \RegFile/_6788_ ( .A(\RegFile/_2687_ ), .B1(\RegFile/_2146_ ), .B2(\RegFile/_2688_ ), .ZN(\RegFile/_2689_ ) );
AOI221_X4 \RegFile/_6789_ ( .A(\RegFile/_2689_ ), .B1(\RegFile/_3657_ ), .B2(\RegFile/_2133_ ), .C1(\RegFile/_3305_ ), .C2(\RegFile/_2066_ ), .ZN(\RegFile/_2690_ ) );
AOI22_X1 \RegFile/_6790_ ( .A1(\RegFile/_2085_ ), .A2(\RegFile/_3433_ ), .B1(\RegFile/_2053_ ), .B2(\RegFile/_3625_ ), .ZN(\RegFile/_2691_ ) );
AOI22_X1 \RegFile/_6791_ ( .A1(\RegFile/_2048_ ), .A2(\RegFile/_3529_ ), .B1(\RegFile/_3401_ ), .B2(\RegFile/_2086_ ), .ZN(\RegFile/_2692_ ) );
NAND3_X1 \RegFile/_6792_ ( .A1(\RegFile/_2268_ ), .A2(\RegFile/_3337_ ), .A3(\RegFile/_2254_ ), .ZN(\RegFile/_2693_ ) );
AND4_X1 \RegFile/_6793_ ( .A1(\RegFile/_2062_ ), .A2(\RegFile/_2691_ ), .A3(\RegFile/_2692_ ), .A4(\RegFile/_2693_ ), .ZN(\RegFile/_2694_ ) );
AND3_X1 \RegFile/_6794_ ( .A1(\RegFile/_2117_ ), .A2(\RegFile/_2106_ ), .A3(\RegFile/_3689_ ), .ZN(\RegFile/_2695_ ) );
AOI221_X4 \RegFile/_6795_ ( .A(\RegFile/_2695_ ), .B1(\RegFile/_2008_ ), .B2(\RegFile/_3721_ ), .C1(\RegFile/_3785_ ), .C2(\RegFile/_2014_ ), .ZN(\RegFile/_2696_ ) );
NAND3_X1 \RegFile/_6796_ ( .A1(\RegFile/_2166_ ), .A2(\RegFile/_2170_ ), .A3(\RegFile/_3497_ ), .ZN(\RegFile/_2697_ ) );
NAND3_X1 \RegFile/_6797_ ( .A1(\RegFile/_2268_ ), .A2(\RegFile/_3753_ ), .A3(\RegFile/_2163_ ), .ZN(\RegFile/_2698_ ) );
NAND3_X1 \RegFile/_6798_ ( .A1(\RegFile/_2268_ ), .A2(\RegFile/_3369_ ), .A3(\RegFile/_1989_ ), .ZN(\RegFile/_2699_ ) );
NAND3_X1 \RegFile/_6799_ ( .A1(\RegFile/_2254_ ), .A2(\RegFile/_3465_ ), .A3(\RegFile/_2255_ ), .ZN(\RegFile/_2700_ ) );
AND4_X1 \RegFile/_6800_ ( .A1(\RegFile/_2697_ ), .A2(\RegFile/_2698_ ), .A3(\RegFile/_2699_ ), .A4(\RegFile/_2700_ ), .ZN(\RegFile/_2701_ ) );
NAND4_X4 \RegFile/_6801_ ( .A1(\RegFile/_2690_ ), .A2(\RegFile/_2694_ ), .A3(\RegFile/_2696_ ), .A4(\RegFile/_2701_ ), .ZN(\RegFile/_2702_ ) );
OR3_X1 \RegFile/_6802_ ( .A1(\RegFile/_2236_ ), .A2(\RegFile/_2237_ ), .A3(\RegFile/_0739_ ), .ZN(\RegFile/_2703_ ) );
NAND2_X4 \RegFile/_6803_ ( .A1(\RegFile/_2702_ ), .A2(\RegFile/_2703_ ), .ZN(\RegFile/_2704_ ) );
BUF_X4 \RegFile/_6804_ ( .A(\RegFile/_2704_ ), .Z(\RegFile/_2705_ ) );
OAI21_X1 \RegFile/_6805_ ( .A(\RegFile/_2686_ ), .B1(\RegFile/_2705_ ), .B2(\RegFile/_2077_ ), .ZN(\RegFile/_0638_ ) );
BUF_X4 \RegFile/_6806_ ( .A(\RegFile/_1990_ ), .Z(\RegFile/_2706_ ) );
AOI21_X1 \RegFile/_6807_ ( .A(\RegFile/_3498_ ), .B1(\RegFile/_2706_ ), .B2(\RegFile/_2665_ ), .ZN(\RegFile/_2707_ ) );
NAND3_X1 \RegFile/_6808_ ( .A1(\RegFile/_2220_ ), .A2(\RegFile/_3626_ ), .A3(\RegFile/_2034_ ), .ZN(\RegFile/_2708_ ) );
OAI21_X1 \RegFile/_6809_ ( .A(\RegFile/_2708_ ), .B1(\RegFile/_2182_ ), .B2(\RegFile/_1378_ ), .ZN(\RegFile/_2709_ ) );
AOI221_X1 \RegFile/_6810_ ( .A(\RegFile/_2709_ ), .B1(\RegFile/_3594_ ), .B2(\RegFile/_2177_ ), .C1(\RegFile/_3562_ ), .C2(\RegFile/_2228_ ), .ZN(\RegFile/_2710_ ) );
AOI22_X1 \RegFile/_6811_ ( .A1(\RegFile/_2155_ ), .A2(\RegFile/_3530_ ), .B1(\RegFile/_3306_ ), .B2(\RegFile/_2121_ ), .ZN(\RegFile/_2711_ ) );
AOI22_X1 \RegFile/_6812_ ( .A1(\RegFile/_3338_ ), .A2(\RegFile/_2018_ ), .B1(\RegFile/_2081_ ), .B2(\RegFile/_3370_ ), .ZN(\RegFile/_2712_ ) );
AND3_X1 \RegFile/_6813_ ( .A1(\RegFile/_2040_ ), .A2(\RegFile/_2041_ ), .A3(\RegFile/_3690_ ), .ZN(\RegFile/_2713_ ) );
AOI21_X1 \RegFile/_6814_ ( .A(\RegFile/_2713_ ), .B1(\RegFile/_3722_ ), .B2(\RegFile/_2009_ ), .ZN(\RegFile/_2714_ ) );
AOI22_X1 \RegFile/_6815_ ( .A1(\RegFile/_2085_ ), .A2(\RegFile/_3434_ ), .B1(\RegFile/_3402_ ), .B2(\RegFile/_2086_ ), .ZN(\RegFile/_2715_ ) );
AND4_X1 \RegFile/_6816_ ( .A1(\RegFile/_2711_ ), .A2(\RegFile/_2712_ ), .A3(\RegFile/_2714_ ), .A4(\RegFile/_2715_ ), .ZN(\RegFile/_2716_ ) );
NAND3_X1 \RegFile/_6817_ ( .A1(\RegFile/_2041_ ), .A2(\RegFile/_3466_ ), .A3(\RegFile/_2103_ ), .ZN(\RegFile/_2717_ ) );
NAND3_X1 \RegFile/_6818_ ( .A1(\RegFile/_1988_ ), .A2(\RegFile/_2103_ ), .A3(\RegFile/_3498_ ), .ZN(\RegFile/_2718_ ) );
NAND2_X1 \RegFile/_6819_ ( .A1(\RegFile/_2717_ ), .A2(\RegFile/_2718_ ), .ZN(\RegFile/_2719_ ) );
AOI221_X4 \RegFile/_6820_ ( .A(\RegFile/_2719_ ), .B1(\RegFile/_2130_ ), .B2(\RegFile/_3786_ ), .C1(\RegFile/_3754_ ), .C2(\RegFile/_2131_ ), .ZN(\RegFile/_2720_ ) );
NAND4_X1 \RegFile/_6821_ ( .A1(\RegFile/_2710_ ), .A2(\RegFile/_2063_ ), .A3(\RegFile/_2716_ ), .A4(\RegFile/_2720_ ), .ZN(\RegFile/_2721_ ) );
OR3_X1 \RegFile/_6822_ ( .A1(\RegFile/_2067_ ), .A2(\RegFile/_2069_ ), .A3(\RegFile/_0740_ ), .ZN(\RegFile/_2722_ ) );
NAND2_X2 \RegFile/_6823_ ( .A1(\RegFile/_2721_ ), .A2(\RegFile/_2722_ ), .ZN(\RegFile/_2723_ ) );
BUF_X4 \RegFile/_6824_ ( .A(\RegFile/_2723_ ), .Z(\RegFile/_2724_ ) );
AOI21_X1 \RegFile/_6825_ ( .A(\RegFile/_2707_ ), .B1(\RegFile/_2724_ ), .B2(\RegFile/_2074_ ), .ZN(\RegFile/_0639_ ) );
CLKBUF_X1 \RegFile/_6826_ ( .A(\RegFile/_3282_ ), .Z(\RegFile/_0128_ ) );
CLKBUF_X1 \RegFile/_6827_ ( .A(\RegFile/_3293_ ), .Z(\RegFile/_0129_ ) );
CLKBUF_X1 \RegFile/_6828_ ( .A(\RegFile/_3304_ ), .Z(\RegFile/_0130_ ) );
CLKBUF_X1 \RegFile/_6829_ ( .A(\RegFile/_3307_ ), .Z(\RegFile/_0131_ ) );
CLKBUF_X1 \RegFile/_6830_ ( .A(\RegFile/_3308_ ), .Z(\RegFile/_0132_ ) );
CLKBUF_X1 \RegFile/_6831_ ( .A(\RegFile/_3309_ ), .Z(\RegFile/_0133_ ) );
CLKBUF_X1 \RegFile/_6832_ ( .A(\RegFile/_3310_ ), .Z(\RegFile/_0134_ ) );
CLKBUF_X1 \RegFile/_6833_ ( .A(\RegFile/_3311_ ), .Z(\RegFile/_0135_ ) );
CLKBUF_X1 \RegFile/_6834_ ( .A(\RegFile/_3312_ ), .Z(\RegFile/_0136_ ) );
CLKBUF_X1 \RegFile/_6835_ ( .A(\RegFile/_3313_ ), .Z(\RegFile/_0137_ ) );
CLKBUF_X1 \RegFile/_6836_ ( .A(\RegFile/_3283_ ), .Z(\RegFile/_0138_ ) );
CLKBUF_X1 \RegFile/_6837_ ( .A(\RegFile/_3284_ ), .Z(\RegFile/_0139_ ) );
CLKBUF_X1 \RegFile/_6838_ ( .A(\RegFile/_3285_ ), .Z(\RegFile/_0140_ ) );
CLKBUF_X1 \RegFile/_6839_ ( .A(\RegFile/_3286_ ), .Z(\RegFile/_0141_ ) );
CLKBUF_X1 \RegFile/_6840_ ( .A(\RegFile/_3287_ ), .Z(\RegFile/_0142_ ) );
CLKBUF_X1 \RegFile/_6841_ ( .A(\RegFile/_3288_ ), .Z(\RegFile/_0143_ ) );
CLKBUF_X1 \RegFile/_6842_ ( .A(\RegFile/_3289_ ), .Z(\RegFile/_0144_ ) );
CLKBUF_X1 \RegFile/_6843_ ( .A(\RegFile/_3290_ ), .Z(\RegFile/_0145_ ) );
CLKBUF_X1 \RegFile/_6844_ ( .A(\RegFile/_3291_ ), .Z(\RegFile/_0146_ ) );
CLKBUF_X1 \RegFile/_6845_ ( .A(\RegFile/_3292_ ), .Z(\RegFile/_0147_ ) );
CLKBUF_X1 \RegFile/_6846_ ( .A(\RegFile/_3294_ ), .Z(\RegFile/_0148_ ) );
CLKBUF_X1 \RegFile/_6847_ ( .A(\RegFile/_3295_ ), .Z(\RegFile/_0149_ ) );
CLKBUF_X1 \RegFile/_6848_ ( .A(\RegFile/_3296_ ), .Z(\RegFile/_0150_ ) );
CLKBUF_X1 \RegFile/_6849_ ( .A(\RegFile/_3297_ ), .Z(\RegFile/_0151_ ) );
CLKBUF_X1 \RegFile/_6850_ ( .A(\RegFile/_3298_ ), .Z(\RegFile/_0152_ ) );
CLKBUF_X1 \RegFile/_6851_ ( .A(\RegFile/_3299_ ), .Z(\RegFile/_0153_ ) );
CLKBUF_X1 \RegFile/_6852_ ( .A(\RegFile/_3300_ ), .Z(\RegFile/_0154_ ) );
CLKBUF_X1 \RegFile/_6853_ ( .A(\RegFile/_3301_ ), .Z(\RegFile/_0155_ ) );
CLKBUF_X1 \RegFile/_6854_ ( .A(\RegFile/_3302_ ), .Z(\RegFile/_0156_ ) );
CLKBUF_X1 \RegFile/_6855_ ( .A(\RegFile/_3303_ ), .Z(\RegFile/_0157_ ) );
CLKBUF_X1 \RegFile/_6856_ ( .A(\RegFile/_3305_ ), .Z(\RegFile/_0158_ ) );
CLKBUF_X1 \RegFile/_6857_ ( .A(\RegFile/_3306_ ), .Z(\RegFile/_0159_ ) );
BUF_X4 \RegFile/_6858_ ( .A(\RegFile/_2161_ ), .Z(\RegFile/_2725_ ) );
BUF_X4 \RegFile/_6859_ ( .A(\RegFile/_2725_ ), .Z(\RegFile/_2726_ ) );
BUF_X4 \RegFile/_6860_ ( .A(\RegFile/_2376_ ), .Z(\RegFile/_2727_ ) );
AOI21_X1 \RegFile/_6861_ ( .A(\RegFile/_3506_ ), .B1(\RegFile/_2726_ ), .B2(\RegFile/_2727_ ), .ZN(\RegFile/_2728_ ) );
BUF_X4 \RegFile/_6862_ ( .A(\RegFile/_2155_ ), .Z(\RegFile/_2729_ ) );
BUF_X4 \RegFile/_6863_ ( .A(\RegFile/_2729_ ), .Z(\RegFile/_2730_ ) );
AOI21_X1 \RegFile/_6864_ ( .A(\RegFile/_2728_ ), .B1(\RegFile/_2072_ ), .B2(\RegFile/_2730_ ), .ZN(\RegFile/_0160_ ) );
AOI21_X1 \RegFile/_6865_ ( .A(\RegFile/_3517_ ), .B1(\RegFile/_2726_ ), .B2(\RegFile/_2727_ ), .ZN(\RegFile/_2731_ ) );
AOI21_X1 \RegFile/_6866_ ( .A(\RegFile/_2731_ ), .B1(\RegFile/_2113_ ), .B2(\RegFile/_2730_ ), .ZN(\RegFile/_0161_ ) );
AOI21_X1 \RegFile/_6867_ ( .A(\RegFile/_3528_ ), .B1(\RegFile/_2726_ ), .B2(\RegFile/_2727_ ), .ZN(\RegFile/_2732_ ) );
AOI21_X1 \RegFile/_6868_ ( .A(\RegFile/_2732_ ), .B1(\RegFile/_2142_ ), .B2(\RegFile/_2730_ ), .ZN(\RegFile/_0162_ ) );
AOI21_X1 \RegFile/_6869_ ( .A(\RegFile/_3531_ ), .B1(\RegFile/_2726_ ), .B2(\RegFile/_2727_ ), .ZN(\RegFile/_2733_ ) );
AOI21_X1 \RegFile/_6870_ ( .A(\RegFile/_2733_ ), .B1(\RegFile/_2175_ ), .B2(\RegFile/_2730_ ), .ZN(\RegFile/_0163_ ) );
INV_X2 \RegFile/_6871_ ( .A(\RegFile/_2155_ ), .ZN(\RegFile/_2734_ ) );
BUF_X4 \RegFile/_6872_ ( .A(\RegFile/_2734_ ), .Z(\RegFile/_2735_ ) );
NAND2_X1 \RegFile/_6873_ ( .A1(\RegFile/_2735_ ), .A2(\RegFile/_3532_ ), .ZN(\RegFile/_2736_ ) );
BUF_X4 \RegFile/_6874_ ( .A(\RegFile/_2734_ ), .Z(\RegFile/_2737_ ) );
OAI21_X1 \RegFile/_6875_ ( .A(\RegFile/_2736_ ), .B1(\RegFile/_2199_ ), .B2(\RegFile/_2737_ ), .ZN(\RegFile/_0164_ ) );
AOI21_X1 \RegFile/_6876_ ( .A(\RegFile/_3533_ ), .B1(\RegFile/_2726_ ), .B2(\RegFile/_2727_ ), .ZN(\RegFile/_2738_ ) );
AOI21_X1 \RegFile/_6877_ ( .A(\RegFile/_2738_ ), .B1(\RegFile/_2218_ ), .B2(\RegFile/_2730_ ), .ZN(\RegFile/_0165_ ) );
AOI21_X1 \RegFile/_6878_ ( .A(\RegFile/_3534_ ), .B1(\RegFile/_2726_ ), .B2(\RegFile/_2727_ ), .ZN(\RegFile/_2739_ ) );
AOI21_X1 \RegFile/_6879_ ( .A(\RegFile/_2739_ ), .B1(\RegFile/_2240_ ), .B2(\RegFile/_2730_ ), .ZN(\RegFile/_0166_ ) );
NAND2_X1 \RegFile/_6880_ ( .A1(\RegFile/_2735_ ), .A2(\RegFile/_3535_ ), .ZN(\RegFile/_2740_ ) );
OAI21_X1 \RegFile/_6881_ ( .A(\RegFile/_2740_ ), .B1(\RegFile/_2260_ ), .B2(\RegFile/_2737_ ), .ZN(\RegFile/_0167_ ) );
NAND2_X1 \RegFile/_6882_ ( .A1(\RegFile/_2735_ ), .A2(\RegFile/_3536_ ), .ZN(\RegFile/_2741_ ) );
OAI21_X1 \RegFile/_6883_ ( .A(\RegFile/_2741_ ), .B1(\RegFile/_2280_ ), .B2(\RegFile/_2737_ ), .ZN(\RegFile/_0168_ ) );
NAND2_X1 \RegFile/_6884_ ( .A1(\RegFile/_2735_ ), .A2(\RegFile/_3537_ ), .ZN(\RegFile/_2742_ ) );
OAI21_X1 \RegFile/_6885_ ( .A(\RegFile/_2742_ ), .B1(\RegFile/_2299_ ), .B2(\RegFile/_2737_ ), .ZN(\RegFile/_0169_ ) );
AOI21_X1 \RegFile/_6886_ ( .A(\RegFile/_3507_ ), .B1(\RegFile/_2726_ ), .B2(\RegFile/_2727_ ), .ZN(\RegFile/_2743_ ) );
AOI21_X1 \RegFile/_6887_ ( .A(\RegFile/_2743_ ), .B1(\RegFile/_2318_ ), .B2(\RegFile/_2730_ ), .ZN(\RegFile/_0170_ ) );
AOI21_X1 \RegFile/_6888_ ( .A(\RegFile/_3508_ ), .B1(\RegFile/_2726_ ), .B2(\RegFile/_2727_ ), .ZN(\RegFile/_2744_ ) );
AOI21_X1 \RegFile/_6889_ ( .A(\RegFile/_2744_ ), .B1(\RegFile/_2336_ ), .B2(\RegFile/_2730_ ), .ZN(\RegFile/_0171_ ) );
NAND2_X1 \RegFile/_6890_ ( .A1(\RegFile/_2735_ ), .A2(\RegFile/_3509_ ), .ZN(\RegFile/_2745_ ) );
OAI21_X1 \RegFile/_6891_ ( .A(\RegFile/_2745_ ), .B1(\RegFile/_2356_ ), .B2(\RegFile/_2737_ ), .ZN(\RegFile/_0172_ ) );
NAND2_X1 \RegFile/_6892_ ( .A1(\RegFile/_2735_ ), .A2(\RegFile/_3510_ ), .ZN(\RegFile/_2746_ ) );
OAI21_X1 \RegFile/_6893_ ( .A(\RegFile/_2746_ ), .B1(\RegFile/_2379_ ), .B2(\RegFile/_2737_ ), .ZN(\RegFile/_0173_ ) );
AOI21_X1 \RegFile/_6894_ ( .A(\RegFile/_3511_ ), .B1(\RegFile/_2726_ ), .B2(\RegFile/_2727_ ), .ZN(\RegFile/_2747_ ) );
AOI21_X1 \RegFile/_6895_ ( .A(\RegFile/_2747_ ), .B1(\RegFile/_2399_ ), .B2(\RegFile/_2730_ ), .ZN(\RegFile/_0174_ ) );
AOI21_X1 \RegFile/_6896_ ( .A(\RegFile/_3512_ ), .B1(\RegFile/_2726_ ), .B2(\RegFile/_2727_ ), .ZN(\RegFile/_2748_ ) );
AOI21_X1 \RegFile/_6897_ ( .A(\RegFile/_2748_ ), .B1(\RegFile/_2420_ ), .B2(\RegFile/_2730_ ), .ZN(\RegFile/_0175_ ) );
BUF_X4 \RegFile/_6898_ ( .A(\RegFile/_2725_ ), .Z(\RegFile/_2749_ ) );
BUF_X4 \RegFile/_6899_ ( .A(\RegFile/_2376_ ), .Z(\RegFile/_2750_ ) );
AOI21_X1 \RegFile/_6900_ ( .A(\RegFile/_3513_ ), .B1(\RegFile/_2749_ ), .B2(\RegFile/_2750_ ), .ZN(\RegFile/_2751_ ) );
AOI21_X1 \RegFile/_6901_ ( .A(\RegFile/_2751_ ), .B1(\RegFile/_2440_ ), .B2(\RegFile/_2729_ ), .ZN(\RegFile/_0176_ ) );
AOI21_X1 \RegFile/_6902_ ( .A(\RegFile/_3514_ ), .B1(\RegFile/_2749_ ), .B2(\RegFile/_2750_ ), .ZN(\RegFile/_2752_ ) );
AOI21_X1 \RegFile/_6903_ ( .A(\RegFile/_2752_ ), .B1(\RegFile/_2459_ ), .B2(\RegFile/_2729_ ), .ZN(\RegFile/_0177_ ) );
AOI21_X1 \RegFile/_6904_ ( .A(\RegFile/_3515_ ), .B1(\RegFile/_2749_ ), .B2(\RegFile/_2750_ ), .ZN(\RegFile/_2753_ ) );
AOI21_X1 \RegFile/_6905_ ( .A(\RegFile/_2753_ ), .B1(\RegFile/_2476_ ), .B2(\RegFile/_2729_ ), .ZN(\RegFile/_0178_ ) );
NAND2_X1 \RegFile/_6906_ ( .A1(\RegFile/_2735_ ), .A2(\RegFile/_3516_ ), .ZN(\RegFile/_2754_ ) );
OAI21_X1 \RegFile/_6907_ ( .A(\RegFile/_2754_ ), .B1(\RegFile/_2495_ ), .B2(\RegFile/_2737_ ), .ZN(\RegFile/_0179_ ) );
NAND2_X1 \RegFile/_6908_ ( .A1(\RegFile/_2734_ ), .A2(\RegFile/_3518_ ), .ZN(\RegFile/_2755_ ) );
OAI21_X1 \RegFile/_6909_ ( .A(\RegFile/_2755_ ), .B1(\RegFile/_2514_ ), .B2(\RegFile/_2737_ ), .ZN(\RegFile/_0180_ ) );
NAND2_X1 \RegFile/_6910_ ( .A1(\RegFile/_2734_ ), .A2(\RegFile/_3519_ ), .ZN(\RegFile/_2756_ ) );
OAI21_X1 \RegFile/_6911_ ( .A(\RegFile/_2756_ ), .B1(\RegFile/_2533_ ), .B2(\RegFile/_2737_ ), .ZN(\RegFile/_0181_ ) );
AOI21_X1 \RegFile/_6912_ ( .A(\RegFile/_3520_ ), .B1(\RegFile/_2749_ ), .B2(\RegFile/_2750_ ), .ZN(\RegFile/_2757_ ) );
AOI21_X1 \RegFile/_6913_ ( .A(\RegFile/_2757_ ), .B1(\RegFile/_2552_ ), .B2(\RegFile/_2729_ ), .ZN(\RegFile/_0182_ ) );
AOI21_X1 \RegFile/_6914_ ( .A(\RegFile/_3521_ ), .B1(\RegFile/_2749_ ), .B2(\RegFile/_2750_ ), .ZN(\RegFile/_2758_ ) );
AOI21_X1 \RegFile/_6915_ ( .A(\RegFile/_2758_ ), .B1(\RegFile/_2571_ ), .B2(\RegFile/_2729_ ), .ZN(\RegFile/_0183_ ) );
NAND2_X1 \RegFile/_6916_ ( .A1(\RegFile/_2734_ ), .A2(\RegFile/_3522_ ), .ZN(\RegFile/_2759_ ) );
OAI21_X1 \RegFile/_6917_ ( .A(\RegFile/_2759_ ), .B1(\RegFile/_2592_ ), .B2(\RegFile/_2737_ ), .ZN(\RegFile/_0184_ ) );
AOI21_X1 \RegFile/_6918_ ( .A(\RegFile/_3523_ ), .B1(\RegFile/_2749_ ), .B2(\RegFile/_2750_ ), .ZN(\RegFile/_2760_ ) );
AOI21_X1 \RegFile/_6919_ ( .A(\RegFile/_2760_ ), .B1(\RegFile/_2608_ ), .B2(\RegFile/_2729_ ), .ZN(\RegFile/_0185_ ) );
NAND2_X1 \RegFile/_6920_ ( .A1(\RegFile/_2734_ ), .A2(\RegFile/_3524_ ), .ZN(\RegFile/_2761_ ) );
OAI21_X1 \RegFile/_6921_ ( .A(\RegFile/_2761_ ), .B1(\RegFile/_2628_ ), .B2(\RegFile/_2735_ ), .ZN(\RegFile/_0186_ ) );
AOI21_X1 \RegFile/_6922_ ( .A(\RegFile/_3525_ ), .B1(\RegFile/_2749_ ), .B2(\RegFile/_2750_ ), .ZN(\RegFile/_2762_ ) );
AOI21_X1 \RegFile/_6923_ ( .A(\RegFile/_2762_ ), .B1(\RegFile/_2646_ ), .B2(\RegFile/_2729_ ), .ZN(\RegFile/_0187_ ) );
AOI21_X1 \RegFile/_6924_ ( .A(\RegFile/_3526_ ), .B1(\RegFile/_2749_ ), .B2(\RegFile/_2750_ ), .ZN(\RegFile/_2763_ ) );
AOI21_X1 \RegFile/_6925_ ( .A(\RegFile/_2763_ ), .B1(\RegFile/_2664_ ), .B2(\RegFile/_2729_ ), .ZN(\RegFile/_0188_ ) );
NAND2_X1 \RegFile/_6926_ ( .A1(\RegFile/_2734_ ), .A2(\RegFile/_3527_ ), .ZN(\RegFile/_2764_ ) );
OAI21_X1 \RegFile/_6927_ ( .A(\RegFile/_2764_ ), .B1(\RegFile/_2685_ ), .B2(\RegFile/_2735_ ), .ZN(\RegFile/_0189_ ) );
NAND2_X1 \RegFile/_6928_ ( .A1(\RegFile/_2734_ ), .A2(\RegFile/_3529_ ), .ZN(\RegFile/_2765_ ) );
OAI21_X1 \RegFile/_6929_ ( .A(\RegFile/_2765_ ), .B1(\RegFile/_2705_ ), .B2(\RegFile/_2735_ ), .ZN(\RegFile/_0190_ ) );
AOI21_X1 \RegFile/_6930_ ( .A(\RegFile/_3530_ ), .B1(\RegFile/_2749_ ), .B2(\RegFile/_2750_ ), .ZN(\RegFile/_2766_ ) );
AOI21_X1 \RegFile/_6931_ ( .A(\RegFile/_2766_ ), .B1(\RegFile/_2724_ ), .B2(\RegFile/_2729_ ), .ZN(\RegFile/_0191_ ) );
BUF_X4 \RegFile/_6932_ ( .A(\RegFile/_2169_ ), .Z(\RegFile/_2767_ ) );
AOI21_X1 \RegFile/_6933_ ( .A(\RegFile/_3538_ ), .B1(\RegFile/_2767_ ), .B2(\RegFile/_2750_ ), .ZN(\RegFile/_2768_ ) );
BUF_X4 \RegFile/_6934_ ( .A(\RegFile/_2228_ ), .Z(\RegFile/_2769_ ) );
AOI21_X1 \RegFile/_6935_ ( .A(\RegFile/_2768_ ), .B1(\RegFile/_2072_ ), .B2(\RegFile/_2769_ ), .ZN(\RegFile/_0192_ ) );
BUF_X4 \RegFile/_6936_ ( .A(\RegFile/_2376_ ), .Z(\RegFile/_2770_ ) );
AOI21_X1 \RegFile/_6937_ ( .A(\RegFile/_3549_ ), .B1(\RegFile/_2767_ ), .B2(\RegFile/_2770_ ), .ZN(\RegFile/_2771_ ) );
AOI21_X1 \RegFile/_6938_ ( .A(\RegFile/_2771_ ), .B1(\RegFile/_2113_ ), .B2(\RegFile/_2769_ ), .ZN(\RegFile/_0193_ ) );
AOI21_X1 \RegFile/_6939_ ( .A(\RegFile/_3560_ ), .B1(\RegFile/_2767_ ), .B2(\RegFile/_2770_ ), .ZN(\RegFile/_2772_ ) );
AOI21_X1 \RegFile/_6940_ ( .A(\RegFile/_2772_ ), .B1(\RegFile/_2142_ ), .B2(\RegFile/_2769_ ), .ZN(\RegFile/_0194_ ) );
BUF_X4 \RegFile/_6941_ ( .A(\RegFile/_2228_ ), .Z(\RegFile/_2773_ ) );
NAND3_X1 \RegFile/_6942_ ( .A1(\RegFile/_2173_ ), .A2(\RegFile/_2773_ ), .A3(\RegFile/_2174_ ), .ZN(\RegFile/_2774_ ) );
OAI21_X1 \RegFile/_6943_ ( .A(\RegFile/_2774_ ), .B1(\RegFile/_1511_ ), .B2(\RegFile/_2773_ ), .ZN(\RegFile/_0195_ ) );
AND2_X1 \RegFile/_6944_ ( .A1(\RegFile/_2198_ ), .A2(\RegFile/_2228_ ), .ZN(\RegFile/_2775_ ) );
BUF_X4 \RegFile/_6945_ ( .A(\RegFile/_2362_ ), .Z(\RegFile/_2776_ ) );
AOI21_X1 \RegFile/_6946_ ( .A(\RegFile/_2775_ ), .B1(\RegFile/_0915_ ), .B2(\RegFile/_2776_ ), .ZN(\RegFile/_0196_ ) );
AOI21_X1 \RegFile/_6947_ ( .A(\RegFile/_2362_ ), .B1(\RegFile/_2216_ ), .B2(\RegFile/_2217_ ), .ZN(\RegFile/_2777_ ) );
AOI21_X1 \RegFile/_6948_ ( .A(\RegFile/_2777_ ), .B1(\RegFile/_1546_ ), .B2(\RegFile/_2776_ ), .ZN(\RegFile/_0197_ ) );
BUF_X4 \RegFile/_6949_ ( .A(\RegFile/_2362_ ), .Z(\RegFile/_2778_ ) );
NAND2_X1 \RegFile/_6950_ ( .A1(\RegFile/_2778_ ), .A2(\RegFile/_3566_ ), .ZN(\RegFile/_2779_ ) );
OAI21_X1 \RegFile/_6951_ ( .A(\RegFile/_2779_ ), .B1(\RegFile/_2240_ ), .B2(\RegFile/_2776_ ), .ZN(\RegFile/_0198_ ) );
AOI21_X1 \RegFile/_6952_ ( .A(\RegFile/_3567_ ), .B1(\RegFile/_2767_ ), .B2(\RegFile/_2770_ ), .ZN(\RegFile/_2780_ ) );
AOI21_X1 \RegFile/_6953_ ( .A(\RegFile/_2780_ ), .B1(\RegFile/_2261_ ), .B2(\RegFile/_2769_ ), .ZN(\RegFile/_0199_ ) );
AOI21_X1 \RegFile/_6954_ ( .A(\RegFile/_3568_ ), .B1(\RegFile/_2767_ ), .B2(\RegFile/_2770_ ), .ZN(\RegFile/_2781_ ) );
BUF_X4 \RegFile/_6955_ ( .A(\RegFile/_2280_ ), .Z(\RegFile/_2782_ ) );
AOI21_X1 \RegFile/_6956_ ( .A(\RegFile/_2781_ ), .B1(\RegFile/_2782_ ), .B2(\RegFile/_2769_ ), .ZN(\RegFile/_0200_ ) );
AOI21_X1 \RegFile/_6957_ ( .A(\RegFile/_3569_ ), .B1(\RegFile/_2767_ ), .B2(\RegFile/_2770_ ), .ZN(\RegFile/_2783_ ) );
AOI21_X1 \RegFile/_6958_ ( .A(\RegFile/_2783_ ), .B1(\RegFile/_2299_ ), .B2(\RegFile/_2769_ ), .ZN(\RegFile/_0201_ ) );
AOI21_X1 \RegFile/_6959_ ( .A(\RegFile/_3539_ ), .B1(\RegFile/_2767_ ), .B2(\RegFile/_2770_ ), .ZN(\RegFile/_2784_ ) );
AOI21_X1 \RegFile/_6960_ ( .A(\RegFile/_2784_ ), .B1(\RegFile/_2318_ ), .B2(\RegFile/_2769_ ), .ZN(\RegFile/_0202_ ) );
OR3_X1 \RegFile/_6961_ ( .A1(\RegFile/_2333_ ), .A2(\RegFile/_2362_ ), .A3(\RegFile/_2334_ ), .ZN(\RegFile/_2785_ ) );
OAI21_X1 \RegFile/_6962_ ( .A(\RegFile/_2785_ ), .B1(\RegFile/_1654_ ), .B2(\RegFile/_2773_ ), .ZN(\RegFile/_0203_ ) );
AOI21_X1 \RegFile/_6963_ ( .A(\RegFile/_2362_ ), .B1(\RegFile/_2354_ ), .B2(\RegFile/_2355_ ), .ZN(\RegFile/_2786_ ) );
AOI21_X1 \RegFile/_6964_ ( .A(\RegFile/_2786_ ), .B1(\RegFile/_1059_ ), .B2(\RegFile/_2776_ ), .ZN(\RegFile/_0204_ ) );
AND2_X1 \RegFile/_6965_ ( .A1(\RegFile/_2378_ ), .A2(\RegFile/_2228_ ), .ZN(\RegFile/_2787_ ) );
AOI21_X1 \RegFile/_6966_ ( .A(\RegFile/_2787_ ), .B1(\RegFile/_2361_ ), .B2(\RegFile/_2776_ ), .ZN(\RegFile/_0205_ ) );
AOI21_X1 \RegFile/_6967_ ( .A(\RegFile/_2362_ ), .B1(\RegFile/_2397_ ), .B2(\RegFile/_2398_ ), .ZN(\RegFile/_2788_ ) );
AOI21_X1 \RegFile/_6968_ ( .A(\RegFile/_2788_ ), .B1(\RegFile/_1701_ ), .B2(\RegFile/_2776_ ), .ZN(\RegFile/_0206_ ) );
AOI21_X1 \RegFile/_6969_ ( .A(\RegFile/_3544_ ), .B1(\RegFile/_2767_ ), .B2(\RegFile/_2770_ ), .ZN(\RegFile/_2789_ ) );
AOI21_X1 \RegFile/_6970_ ( .A(\RegFile/_2789_ ), .B1(\RegFile/_2420_ ), .B2(\RegFile/_2769_ ), .ZN(\RegFile/_0207_ ) );
NAND2_X1 \RegFile/_6971_ ( .A1(\RegFile/_2778_ ), .A2(\RegFile/_3545_ ), .ZN(\RegFile/_2790_ ) );
OAI21_X1 \RegFile/_6972_ ( .A(\RegFile/_2790_ ), .B1(\RegFile/_2440_ ), .B2(\RegFile/_2776_ ), .ZN(\RegFile/_0208_ ) );
NAND2_X1 \RegFile/_6973_ ( .A1(\RegFile/_2778_ ), .A2(\RegFile/_3546_ ), .ZN(\RegFile/_2791_ ) );
OAI21_X1 \RegFile/_6974_ ( .A(\RegFile/_2791_ ), .B1(\RegFile/_2459_ ), .B2(\RegFile/_2778_ ), .ZN(\RegFile/_0209_ ) );
AOI21_X1 \RegFile/_6975_ ( .A(\RegFile/_3547_ ), .B1(\RegFile/_2767_ ), .B2(\RegFile/_2770_ ), .ZN(\RegFile/_2792_ ) );
AOI21_X1 \RegFile/_6976_ ( .A(\RegFile/_2792_ ), .B1(\RegFile/_2476_ ), .B2(\RegFile/_2769_ ), .ZN(\RegFile/_0210_ ) );
NAND2_X1 \RegFile/_6977_ ( .A1(\RegFile/_2778_ ), .A2(\RegFile/_3548_ ), .ZN(\RegFile/_2793_ ) );
OAI21_X1 \RegFile/_6978_ ( .A(\RegFile/_2793_ ), .B1(\RegFile/_2495_ ), .B2(\RegFile/_2778_ ), .ZN(\RegFile/_0211_ ) );
AND2_X1 \RegFile/_6979_ ( .A1(\RegFile/_2513_ ), .A2(\RegFile/_2228_ ), .ZN(\RegFile/_2794_ ) );
AOI21_X1 \RegFile/_6980_ ( .A(\RegFile/_2794_ ), .B1(\RegFile/_1807_ ), .B2(\RegFile/_2776_ ), .ZN(\RegFile/_0212_ ) );
AOI21_X1 \RegFile/_6981_ ( .A(\RegFile/_2362_ ), .B1(\RegFile/_2530_ ), .B2(\RegFile/_2531_ ), .ZN(\RegFile/_2795_ ) );
AOI21_X1 \RegFile/_6982_ ( .A(\RegFile/_2795_ ), .B1(\RegFile/_1816_ ), .B2(\RegFile/_2776_ ), .ZN(\RegFile/_0213_ ) );
NAND2_X1 \RegFile/_6983_ ( .A1(\RegFile/_2778_ ), .A2(\RegFile/_3552_ ), .ZN(\RegFile/_2796_ ) );
OAI21_X1 \RegFile/_6984_ ( .A(\RegFile/_2796_ ), .B1(\RegFile/_2552_ ), .B2(\RegFile/_2778_ ), .ZN(\RegFile/_0214_ ) );
NAND3_X1 \RegFile/_6985_ ( .A1(\RegFile/_2568_ ), .A2(\RegFile/_2773_ ), .A3(\RegFile/_2569_ ), .ZN(\RegFile/_2797_ ) );
OAI21_X1 \RegFile/_6986_ ( .A(\RegFile/_2797_ ), .B1(\RegFile/_1854_ ), .B2(\RegFile/_2773_ ), .ZN(\RegFile/_0215_ ) );
AOI21_X1 \RegFile/_6987_ ( .A(\RegFile/_3554_ ), .B1(\RegFile/_2767_ ), .B2(\RegFile/_2770_ ), .ZN(\RegFile/_2798_ ) );
AOI21_X1 \RegFile/_6988_ ( .A(\RegFile/_2798_ ), .B1(\RegFile/_2592_ ), .B2(\RegFile/_2769_ ), .ZN(\RegFile/_0216_ ) );
AOI21_X1 \RegFile/_6989_ ( .A(\RegFile/_2362_ ), .B1(\RegFile/_2606_ ), .B2(\RegFile/_2607_ ), .ZN(\RegFile/_2799_ ) );
AOI21_X1 \RegFile/_6990_ ( .A(\RegFile/_2799_ ), .B1(\RegFile/_1272_ ), .B2(\RegFile/_2776_ ), .ZN(\RegFile/_0217_ ) );
NAND2_X1 \RegFile/_6991_ ( .A1(\RegFile/_2778_ ), .A2(\RegFile/_3556_ ), .ZN(\RegFile/_2800_ ) );
OAI21_X1 \RegFile/_6992_ ( .A(\RegFile/_2800_ ), .B1(\RegFile/_2628_ ), .B2(\RegFile/_2778_ ), .ZN(\RegFile/_0218_ ) );
NAND3_X1 \RegFile/_6993_ ( .A1(\RegFile/_2643_ ), .A2(\RegFile/_2228_ ), .A3(\RegFile/_2644_ ), .ZN(\RegFile/_2801_ ) );
OAI21_X1 \RegFile/_6994_ ( .A(\RegFile/_2801_ ), .B1(\RegFile/_1913_ ), .B2(\RegFile/_2773_ ), .ZN(\RegFile/_0219_ ) );
BUF_X4 \RegFile/_6995_ ( .A(\RegFile/_2169_ ), .Z(\RegFile/_2802_ ) );
AOI21_X1 \RegFile/_6996_ ( .A(\RegFile/_3558_ ), .B1(\RegFile/_2802_ ), .B2(\RegFile/_2770_ ), .ZN(\RegFile/_2803_ ) );
AOI21_X1 \RegFile/_6997_ ( .A(\RegFile/_2803_ ), .B1(\RegFile/_2664_ ), .B2(\RegFile/_2773_ ), .ZN(\RegFile/_0220_ ) );
OR3_X1 \RegFile/_6998_ ( .A1(\RegFile/_2682_ ), .A2(\RegFile/_2362_ ), .A3(\RegFile/_2683_ ), .ZN(\RegFile/_2804_ ) );
OAI21_X1 \RegFile/_6999_ ( .A(\RegFile/_2804_ ), .B1(\RegFile/_2669_ ), .B2(\RegFile/_2773_ ), .ZN(\RegFile/_0221_ ) );
BUF_X4 \RegFile/_7000_ ( .A(\RegFile/_2376_ ), .Z(\RegFile/_2805_ ) );
AOI21_X1 \RegFile/_7001_ ( .A(\RegFile/_3561_ ), .B1(\RegFile/_2802_ ), .B2(\RegFile/_2805_ ), .ZN(\RegFile/_2806_ ) );
AOI21_X1 \RegFile/_7002_ ( .A(\RegFile/_2806_ ), .B1(\RegFile/_2705_ ), .B2(\RegFile/_2773_ ), .ZN(\RegFile/_0222_ ) );
AOI21_X1 \RegFile/_7003_ ( .A(\RegFile/_3562_ ), .B1(\RegFile/_2802_ ), .B2(\RegFile/_2805_ ), .ZN(\RegFile/_2807_ ) );
AOI21_X1 \RegFile/_7004_ ( .A(\RegFile/_2807_ ), .B1(\RegFile/_2724_ ), .B2(\RegFile/_2773_ ), .ZN(\RegFile/_0223_ ) );
AOI21_X1 \RegFile/_7005_ ( .A(\RegFile/_3570_ ), .B1(\RegFile/_2706_ ), .B2(\RegFile/_2805_ ), .ZN(\RegFile/_2808_ ) );
BUF_X4 \RegFile/_7006_ ( .A(\RegFile/_2055_ ), .Z(\RegFile/_2809_ ) );
AOI21_X1 \RegFile/_7007_ ( .A(\RegFile/_2808_ ), .B1(\RegFile/_2072_ ), .B2(\RegFile/_2809_ ), .ZN(\RegFile/_0224_ ) );
BUF_X4 \RegFile/_7008_ ( .A(\RegFile/_2055_ ), .Z(\RegFile/_2810_ ) );
NAND3_X1 \RegFile/_7009_ ( .A1(\RegFile/_2110_ ), .A2(\RegFile/_2810_ ), .A3(\RegFile/_2111_ ), .ZN(\RegFile/_2811_ ) );
BUF_X4 \RegFile/_7010_ ( .A(\RegFile/_2055_ ), .Z(\RegFile/_2812_ ) );
OAI21_X1 \RegFile/_7011_ ( .A(\RegFile/_2811_ ), .B1(\RegFile/_0839_ ), .B2(\RegFile/_2812_ ), .ZN(\RegFile/_0225_ ) );
NAND3_X1 \RegFile/_7012_ ( .A1(\RegFile/_2139_ ), .A2(\RegFile/_2810_ ), .A3(\RegFile/_2140_ ), .ZN(\RegFile/_2813_ ) );
OAI21_X1 \RegFile/_7013_ ( .A(\RegFile/_2813_ ), .B1(\RegFile/_1475_ ), .B2(\RegFile/_2812_ ), .ZN(\RegFile/_0226_ ) );
NAND3_X1 \RegFile/_7014_ ( .A1(\RegFile/_2173_ ), .A2(\RegFile/_2810_ ), .A3(\RegFile/_2174_ ), .ZN(\RegFile/_2814_ ) );
OAI21_X1 \RegFile/_7015_ ( .A(\RegFile/_2814_ ), .B1(\RegFile/_2147_ ), .B2(\RegFile/_2812_ ), .ZN(\RegFile/_0227_ ) );
AOI21_X1 \RegFile/_7016_ ( .A(\RegFile/_3596_ ), .B1(\RegFile/_2706_ ), .B2(\RegFile/_2805_ ), .ZN(\RegFile/_2815_ ) );
AOI21_X1 \RegFile/_7017_ ( .A(\RegFile/_2815_ ), .B1(\RegFile/_2199_ ), .B2(\RegFile/_2809_ ), .ZN(\RegFile/_0228_ ) );
BUF_X4 \RegFile/_7018_ ( .A(\RegFile/_2146_ ), .Z(\RegFile/_2816_ ) );
AOI21_X1 \RegFile/_7019_ ( .A(\RegFile/_2816_ ), .B1(\RegFile/_2216_ ), .B2(\RegFile/_2217_ ), .ZN(\RegFile/_2817_ ) );
BUF_X4 \RegFile/_7020_ ( .A(\RegFile/_2816_ ), .Z(\RegFile/_2818_ ) );
AOI21_X1 \RegFile/_7021_ ( .A(\RegFile/_2817_ ), .B1(\RegFile/_2201_ ), .B2(\RegFile/_2818_ ), .ZN(\RegFile/_0229_ ) );
NAND3_X1 \RegFile/_7022_ ( .A1(\RegFile/_2235_ ), .A2(\RegFile/_2810_ ), .A3(\RegFile/_2238_ ), .ZN(\RegFile/_2819_ ) );
OAI21_X1 \RegFile/_7023_ ( .A(\RegFile/_2819_ ), .B1(\RegFile/_1569_ ), .B2(\RegFile/_2812_ ), .ZN(\RegFile/_0230_ ) );
NAND2_X1 \RegFile/_7024_ ( .A1(\RegFile/_2816_ ), .A2(\RegFile/_3599_ ), .ZN(\RegFile/_2820_ ) );
OAI21_X1 \RegFile/_7025_ ( .A(\RegFile/_2820_ ), .B1(\RegFile/_2260_ ), .B2(\RegFile/_2818_ ), .ZN(\RegFile/_0231_ ) );
AOI21_X1 \RegFile/_7026_ ( .A(\RegFile/_3600_ ), .B1(\RegFile/_2706_ ), .B2(\RegFile/_2805_ ), .ZN(\RegFile/_2821_ ) );
AOI21_X1 \RegFile/_7027_ ( .A(\RegFile/_2821_ ), .B1(\RegFile/_2782_ ), .B2(\RegFile/_2809_ ), .ZN(\RegFile/_0232_ ) );
AOI21_X1 \RegFile/_7028_ ( .A(\RegFile/_3601_ ), .B1(\RegFile/_2706_ ), .B2(\RegFile/_2805_ ), .ZN(\RegFile/_2822_ ) );
AOI21_X1 \RegFile/_7029_ ( .A(\RegFile/_2822_ ), .B1(\RegFile/_2299_ ), .B2(\RegFile/_2809_ ), .ZN(\RegFile/_0233_ ) );
AOI21_X1 \RegFile/_7030_ ( .A(\RegFile/_3571_ ), .B1(\RegFile/_2706_ ), .B2(\RegFile/_2805_ ), .ZN(\RegFile/_2823_ ) );
AOI21_X1 \RegFile/_7031_ ( .A(\RegFile/_2823_ ), .B1(\RegFile/_2318_ ), .B2(\RegFile/_2809_ ), .ZN(\RegFile/_0234_ ) );
AOI21_X1 \RegFile/_7032_ ( .A(\RegFile/_3572_ ), .B1(\RegFile/_2706_ ), .B2(\RegFile/_2805_ ), .ZN(\RegFile/_2824_ ) );
AOI21_X1 \RegFile/_7033_ ( .A(\RegFile/_2824_ ), .B1(\RegFile/_2336_ ), .B2(\RegFile/_2809_ ), .ZN(\RegFile/_0235_ ) );
NAND2_X1 \RegFile/_7034_ ( .A1(\RegFile/_2816_ ), .A2(\RegFile/_3573_ ), .ZN(\RegFile/_2825_ ) );
OAI21_X1 \RegFile/_7035_ ( .A(\RegFile/_2825_ ), .B1(\RegFile/_2356_ ), .B2(\RegFile/_2818_ ), .ZN(\RegFile/_0236_ ) );
AND2_X1 \RegFile/_7036_ ( .A1(\RegFile/_2378_ ), .A2(\RegFile/_2055_ ), .ZN(\RegFile/_2826_ ) );
AOI21_X1 \RegFile/_7037_ ( .A(\RegFile/_2826_ ), .B1(\RegFile/_2360_ ), .B2(\RegFile/_2818_ ), .ZN(\RegFile/_0237_ ) );
NAND3_X1 \RegFile/_7038_ ( .A1(\RegFile/_2397_ ), .A2(\RegFile/_2810_ ), .A3(\RegFile/_2398_ ), .ZN(\RegFile/_2827_ ) );
OAI21_X1 \RegFile/_7039_ ( .A(\RegFile/_2827_ ), .B1(\RegFile/_2390_ ), .B2(\RegFile/_2812_ ), .ZN(\RegFile/_0238_ ) );
NAND2_X1 \RegFile/_7040_ ( .A1(\RegFile/_2816_ ), .A2(\RegFile/_3576_ ), .ZN(\RegFile/_2828_ ) );
OAI21_X1 \RegFile/_7041_ ( .A(\RegFile/_2828_ ), .B1(\RegFile/_2420_ ), .B2(\RegFile/_2818_ ), .ZN(\RegFile/_0239_ ) );
AOI21_X1 \RegFile/_7042_ ( .A(\RegFile/_3577_ ), .B1(\RegFile/_2706_ ), .B2(\RegFile/_2805_ ), .ZN(\RegFile/_2829_ ) );
AOI21_X1 \RegFile/_7043_ ( .A(\RegFile/_2829_ ), .B1(\RegFile/_2440_ ), .B2(\RegFile/_2809_ ), .ZN(\RegFile/_0240_ ) );
OR3_X1 \RegFile/_7044_ ( .A1(\RegFile/_2456_ ), .A2(\RegFile/_2816_ ), .A3(\RegFile/_2457_ ), .ZN(\RegFile/_2830_ ) );
OAI21_X1 \RegFile/_7045_ ( .A(\RegFile/_2830_ ), .B1(\RegFile/_1135_ ), .B2(\RegFile/_2812_ ), .ZN(\RegFile/_0241_ ) );
NAND3_X1 \RegFile/_7046_ ( .A1(\RegFile/_2473_ ), .A2(\RegFile/_2810_ ), .A3(\RegFile/_2474_ ), .ZN(\RegFile/_2831_ ) );
OAI21_X1 \RegFile/_7047_ ( .A(\RegFile/_2831_ ), .B1(\RegFile/_1764_ ), .B2(\RegFile/_2812_ ), .ZN(\RegFile/_0242_ ) );
AND2_X1 \RegFile/_7048_ ( .A1(\RegFile/_2494_ ), .A2(\RegFile/_2055_ ), .ZN(\RegFile/_2832_ ) );
AOI21_X1 \RegFile/_7049_ ( .A(\RegFile/_2832_ ), .B1(\RegFile/_1174_ ), .B2(\RegFile/_2818_ ), .ZN(\RegFile/_0243_ ) );
AOI21_X1 \RegFile/_7050_ ( .A(\RegFile/_3582_ ), .B1(\RegFile/_2706_ ), .B2(\RegFile/_2805_ ), .ZN(\RegFile/_2833_ ) );
AOI21_X1 \RegFile/_7051_ ( .A(\RegFile/_2833_ ), .B1(\RegFile/_2514_ ), .B2(\RegFile/_2809_ ), .ZN(\RegFile/_0244_ ) );
NAND3_X1 \RegFile/_7052_ ( .A1(\RegFile/_2530_ ), .A2(\RegFile/_2810_ ), .A3(\RegFile/_2531_ ), .ZN(\RegFile/_2834_ ) );
OAI21_X1 \RegFile/_7053_ ( .A(\RegFile/_2834_ ), .B1(\RegFile/_2517_ ), .B2(\RegFile/_2812_ ), .ZN(\RegFile/_0245_ ) );
AOI21_X1 \RegFile/_7054_ ( .A(\RegFile/_2816_ ), .B1(\RegFile/_2549_ ), .B2(\RegFile/_2550_ ), .ZN(\RegFile/_2835_ ) );
AOI21_X1 \RegFile/_7055_ ( .A(\RegFile/_2835_ ), .B1(\RegFile/_1833_ ), .B2(\RegFile/_2818_ ), .ZN(\RegFile/_0246_ ) );
AOI21_X1 \RegFile/_7056_ ( .A(\RegFile/_2816_ ), .B1(\RegFile/_2568_ ), .B2(\RegFile/_2569_ ), .ZN(\RegFile/_2836_ ) );
AOI21_X1 \RegFile/_7057_ ( .A(\RegFile/_2836_ ), .B1(\RegFile/_1853_ ), .B2(\RegFile/_2818_ ), .ZN(\RegFile/_0247_ ) );
AOI21_X1 \RegFile/_7058_ ( .A(\RegFile/_3586_ ), .B1(\RegFile/_2706_ ), .B2(\RegFile/_2376_ ), .ZN(\RegFile/_2837_ ) );
AOI21_X1 \RegFile/_7059_ ( .A(\RegFile/_2837_ ), .B1(\RegFile/_2592_ ), .B2(\RegFile/_2809_ ), .ZN(\RegFile/_0248_ ) );
NAND3_X1 \RegFile/_7060_ ( .A1(\RegFile/_2606_ ), .A2(\RegFile/_2810_ ), .A3(\RegFile/_2607_ ), .ZN(\RegFile/_2838_ ) );
OAI21_X1 \RegFile/_7061_ ( .A(\RegFile/_2838_ ), .B1(\RegFile/_1271_ ), .B2(\RegFile/_2810_ ), .ZN(\RegFile/_0249_ ) );
BUF_X4 \RegFile/_7062_ ( .A(\RegFile/_1990_ ), .Z(\RegFile/_2839_ ) );
AOI21_X1 \RegFile/_7063_ ( .A(\RegFile/_3588_ ), .B1(\RegFile/_2839_ ), .B2(\RegFile/_2376_ ), .ZN(\RegFile/_2840_ ) );
AOI21_X1 \RegFile/_7064_ ( .A(\RegFile/_2840_ ), .B1(\RegFile/_2628_ ), .B2(\RegFile/_2809_ ), .ZN(\RegFile/_0250_ ) );
AOI21_X1 \RegFile/_7065_ ( .A(\RegFile/_2816_ ), .B1(\RegFile/_2643_ ), .B2(\RegFile/_2644_ ), .ZN(\RegFile/_2841_ ) );
AOI21_X1 \RegFile/_7066_ ( .A(\RegFile/_2841_ ), .B1(\RegFile/_1912_ ), .B2(\RegFile/_2818_ ), .ZN(\RegFile/_0251_ ) );
AOI21_X1 \RegFile/_7067_ ( .A(\RegFile/_3590_ ), .B1(\RegFile/_2839_ ), .B2(\RegFile/_2376_ ), .ZN(\RegFile/_2842_ ) );
AOI21_X1 \RegFile/_7068_ ( .A(\RegFile/_2842_ ), .B1(\RegFile/_2664_ ), .B2(\RegFile/_2812_ ), .ZN(\RegFile/_0252_ ) );
OR3_X1 \RegFile/_7069_ ( .A1(\RegFile/_2682_ ), .A2(\RegFile/_2146_ ), .A3(\RegFile/_2683_ ), .ZN(\RegFile/_2843_ ) );
OAI21_X1 \RegFile/_7070_ ( .A(\RegFile/_2843_ ), .B1(\RegFile/_2668_ ), .B2(\RegFile/_2810_ ), .ZN(\RegFile/_0253_ ) );
AOI21_X1 \RegFile/_7071_ ( .A(\RegFile/_2816_ ), .B1(\RegFile/_2702_ ), .B2(\RegFile/_2703_ ), .ZN(\RegFile/_2844_ ) );
AOI21_X1 \RegFile/_7072_ ( .A(\RegFile/_2844_ ), .B1(\RegFile/_2688_ ), .B2(\RegFile/_2818_ ), .ZN(\RegFile/_0254_ ) );
AOI21_X1 \RegFile/_7073_ ( .A(\RegFile/_3594_ ), .B1(\RegFile/_2839_ ), .B2(\RegFile/_2376_ ), .ZN(\RegFile/_2845_ ) );
AOI21_X1 \RegFile/_7074_ ( .A(\RegFile/_2845_ ), .B1(\RegFile/_2724_ ), .B2(\RegFile/_2812_ ), .ZN(\RegFile/_0255_ ) );
BUF_X4 \RegFile/_7075_ ( .A(\RegFile/_2338_ ), .Z(\RegFile/_2846_ ) );
BUF_X4 \RegFile/_7076_ ( .A(\RegFile/_2035_ ), .Z(\RegFile/_2847_ ) );
BUF_X4 \RegFile/_7077_ ( .A(\RegFile/_2847_ ), .Z(\RegFile/_2848_ ) );
AOI21_X1 \RegFile/_7078_ ( .A(\RegFile/_3602_ ), .B1(\RegFile/_2846_ ), .B2(\RegFile/_2848_ ), .ZN(\RegFile/_2849_ ) );
BUF_X4 \RegFile/_7079_ ( .A(\RegFile/_2149_ ), .Z(\RegFile/_2850_ ) );
AOI21_X1 \RegFile/_7080_ ( .A(\RegFile/_2849_ ), .B1(\RegFile/_2072_ ), .B2(\RegFile/_2850_ ), .ZN(\RegFile/_0256_ ) );
AOI21_X1 \RegFile/_7081_ ( .A(\RegFile/_3613_ ), .B1(\RegFile/_2846_ ), .B2(\RegFile/_2848_ ), .ZN(\RegFile/_2851_ ) );
AOI21_X1 \RegFile/_7082_ ( .A(\RegFile/_2851_ ), .B1(\RegFile/_2113_ ), .B2(\RegFile/_2850_ ), .ZN(\RegFile/_0257_ ) );
BUF_X4 \RegFile/_7083_ ( .A(\RegFile/_2149_ ), .Z(\RegFile/_2852_ ) );
NAND3_X1 \RegFile/_7084_ ( .A1(\RegFile/_2139_ ), .A2(\RegFile/_2852_ ), .A3(\RegFile/_2140_ ), .ZN(\RegFile/_2853_ ) );
OAI21_X1 \RegFile/_7085_ ( .A(\RegFile/_2853_ ), .B1(\RegFile/_1478_ ), .B2(\RegFile/_2852_ ), .ZN(\RegFile/_0258_ ) );
NAND3_X1 \RegFile/_7086_ ( .A1(\RegFile/_2173_ ), .A2(\RegFile/_2149_ ), .A3(\RegFile/_2174_ ), .ZN(\RegFile/_2854_ ) );
OAI21_X1 \RegFile/_7087_ ( .A(\RegFile/_2854_ ), .B1(\RegFile/_1510_ ), .B2(\RegFile/_2852_ ), .ZN(\RegFile/_0259_ ) );
OR3_X1 \RegFile/_7088_ ( .A1(\RegFile/_2196_ ), .A2(\RegFile/_2180_ ), .A3(\RegFile/_2197_ ), .ZN(\RegFile/_2855_ ) );
OAI21_X1 \RegFile/_7089_ ( .A(\RegFile/_2855_ ), .B1(\RegFile/_0910_ ), .B2(\RegFile/_2852_ ), .ZN(\RegFile/_0260_ ) );
BUF_X4 \RegFile/_7090_ ( .A(\RegFile/_2180_ ), .Z(\RegFile/_2856_ ) );
AOI21_X1 \RegFile/_7091_ ( .A(\RegFile/_2856_ ), .B1(\RegFile/_2216_ ), .B2(\RegFile/_2217_ ), .ZN(\RegFile/_2857_ ) );
BUF_X4 \RegFile/_7092_ ( .A(\RegFile/_2856_ ), .Z(\RegFile/_2858_ ) );
AOI21_X1 \RegFile/_7093_ ( .A(\RegFile/_2857_ ), .B1(\RegFile/_1545_ ), .B2(\RegFile/_2858_ ), .ZN(\RegFile/_0261_ ) );
AOI21_X1 \RegFile/_7094_ ( .A(\RegFile/_2856_ ), .B1(\RegFile/_2235_ ), .B2(\RegFile/_2238_ ), .ZN(\RegFile/_2859_ ) );
AOI21_X1 \RegFile/_7095_ ( .A(\RegFile/_2859_ ), .B1(\RegFile/_1570_ ), .B2(\RegFile/_2858_ ), .ZN(\RegFile/_0262_ ) );
AOI21_X1 \RegFile/_7096_ ( .A(\RegFile/_3631_ ), .B1(\RegFile/_2846_ ), .B2(\RegFile/_2848_ ), .ZN(\RegFile/_2860_ ) );
AOI21_X1 \RegFile/_7097_ ( .A(\RegFile/_2860_ ), .B1(\RegFile/_2261_ ), .B2(\RegFile/_2850_ ), .ZN(\RegFile/_0263_ ) );
AOI21_X1 \RegFile/_7098_ ( .A(\RegFile/_3632_ ), .B1(\RegFile/_2846_ ), .B2(\RegFile/_2848_ ), .ZN(\RegFile/_2861_ ) );
AOI21_X1 \RegFile/_7099_ ( .A(\RegFile/_2861_ ), .B1(\RegFile/_2782_ ), .B2(\RegFile/_2850_ ), .ZN(\RegFile/_0264_ ) );
AOI21_X1 \RegFile/_7100_ ( .A(\RegFile/_2180_ ), .B1(\RegFile/_2296_ ), .B2(\RegFile/_2297_ ), .ZN(\RegFile/_2862_ ) );
AOI21_X1 \RegFile/_7101_ ( .A(\RegFile/_2862_ ), .B1(\RegFile/_1004_ ), .B2(\RegFile/_2858_ ), .ZN(\RegFile/_0265_ ) );
AOI21_X1 \RegFile/_7102_ ( .A(\RegFile/_3603_ ), .B1(\RegFile/_2846_ ), .B2(\RegFile/_2848_ ), .ZN(\RegFile/_2863_ ) );
AOI21_X1 \RegFile/_7103_ ( .A(\RegFile/_2863_ ), .B1(\RegFile/_2318_ ), .B2(\RegFile/_2850_ ), .ZN(\RegFile/_0266_ ) );
AND2_X1 \RegFile/_7104_ ( .A1(\RegFile/_2335_ ), .A2(\RegFile/_2149_ ), .ZN(\RegFile/_2864_ ) );
AOI21_X1 \RegFile/_7105_ ( .A(\RegFile/_2864_ ), .B1(\RegFile/_1653_ ), .B2(\RegFile/_2858_ ), .ZN(\RegFile/_0267_ ) );
AOI21_X1 \RegFile/_7106_ ( .A(\RegFile/_2180_ ), .B1(\RegFile/_2354_ ), .B2(\RegFile/_2355_ ), .ZN(\RegFile/_2865_ ) );
AOI21_X1 \RegFile/_7107_ ( .A(\RegFile/_2865_ ), .B1(\RegFile/_1056_ ), .B2(\RegFile/_2858_ ), .ZN(\RegFile/_0268_ ) );
AOI21_X1 \RegFile/_7108_ ( .A(\RegFile/_3606_ ), .B1(\RegFile/_2846_ ), .B2(\RegFile/_2848_ ), .ZN(\RegFile/_2866_ ) );
AOI21_X1 \RegFile/_7109_ ( .A(\RegFile/_2866_ ), .B1(\RegFile/_2379_ ), .B2(\RegFile/_2850_ ), .ZN(\RegFile/_0269_ ) );
AOI21_X1 \RegFile/_7110_ ( .A(\RegFile/_2180_ ), .B1(\RegFile/_2397_ ), .B2(\RegFile/_2398_ ), .ZN(\RegFile/_2867_ ) );
AOI21_X1 \RegFile/_7111_ ( .A(\RegFile/_2867_ ), .B1(\RegFile/_1700_ ), .B2(\RegFile/_2858_ ), .ZN(\RegFile/_0270_ ) );
AOI21_X1 \RegFile/_7112_ ( .A(\RegFile/_3608_ ), .B1(\RegFile/_2846_ ), .B2(\RegFile/_2848_ ), .ZN(\RegFile/_2868_ ) );
AOI21_X1 \RegFile/_7113_ ( .A(\RegFile/_2868_ ), .B1(\RegFile/_2420_ ), .B2(\RegFile/_2850_ ), .ZN(\RegFile/_0271_ ) );
NAND2_X1 \RegFile/_7114_ ( .A1(\RegFile/_2856_ ), .A2(\RegFile/_3609_ ), .ZN(\RegFile/_2869_ ) );
OAI21_X1 \RegFile/_7115_ ( .A(\RegFile/_2869_ ), .B1(\RegFile/_2440_ ), .B2(\RegFile/_2858_ ), .ZN(\RegFile/_0272_ ) );
AND2_X1 \RegFile/_7116_ ( .A1(\RegFile/_2458_ ), .A2(\RegFile/_2149_ ), .ZN(\RegFile/_2870_ ) );
AOI21_X1 \RegFile/_7117_ ( .A(\RegFile/_2870_ ), .B1(\RegFile/_1136_ ), .B2(\RegFile/_2858_ ), .ZN(\RegFile/_0273_ ) );
AOI21_X1 \RegFile/_7118_ ( .A(\RegFile/_2180_ ), .B1(\RegFile/_2473_ ), .B2(\RegFile/_2474_ ), .ZN(\RegFile/_2871_ ) );
AOI21_X1 \RegFile/_7119_ ( .A(\RegFile/_2871_ ), .B1(\RegFile/_1765_ ), .B2(\RegFile/_2858_ ), .ZN(\RegFile/_0274_ ) );
OR3_X1 \RegFile/_7120_ ( .A1(\RegFile/_2492_ ), .A2(\RegFile/_2180_ ), .A3(\RegFile/_2493_ ), .ZN(\RegFile/_2872_ ) );
OAI21_X1 \RegFile/_7121_ ( .A(\RegFile/_2872_ ), .B1(\RegFile/_1175_ ), .B2(\RegFile/_2852_ ), .ZN(\RegFile/_0275_ ) );
OR3_X1 \RegFile/_7122_ ( .A1(\RegFile/_2511_ ), .A2(\RegFile/_2180_ ), .A3(\RegFile/_2512_ ), .ZN(\RegFile/_2873_ ) );
OAI21_X1 \RegFile/_7123_ ( .A(\RegFile/_2873_ ), .B1(\RegFile/_1806_ ), .B2(\RegFile/_2852_ ), .ZN(\RegFile/_0276_ ) );
NAND3_X1 \RegFile/_7124_ ( .A1(\RegFile/_2530_ ), .A2(\RegFile/_2149_ ), .A3(\RegFile/_2531_ ), .ZN(\RegFile/_2874_ ) );
OAI21_X1 \RegFile/_7125_ ( .A(\RegFile/_2874_ ), .B1(\RegFile/_1815_ ), .B2(\RegFile/_2852_ ), .ZN(\RegFile/_0277_ ) );
AOI21_X1 \RegFile/_7126_ ( .A(\RegFile/_2180_ ), .B1(\RegFile/_2549_ ), .B2(\RegFile/_2550_ ), .ZN(\RegFile/_2875_ ) );
AOI21_X1 \RegFile/_7127_ ( .A(\RegFile/_2875_ ), .B1(\RegFile/_1834_ ), .B2(\RegFile/_2858_ ), .ZN(\RegFile/_0278_ ) );
NAND2_X1 \RegFile/_7128_ ( .A1(\RegFile/_2856_ ), .A2(\RegFile/_3617_ ), .ZN(\RegFile/_2876_ ) );
OAI21_X1 \RegFile/_7129_ ( .A(\RegFile/_2876_ ), .B1(\RegFile/_2571_ ), .B2(\RegFile/_2856_ ), .ZN(\RegFile/_0279_ ) );
NAND2_X1 \RegFile/_7130_ ( .A1(\RegFile/_2856_ ), .A2(\RegFile/_3618_ ), .ZN(\RegFile/_2877_ ) );
OAI21_X1 \RegFile/_7131_ ( .A(\RegFile/_2877_ ), .B1(\RegFile/_2592_ ), .B2(\RegFile/_2856_ ), .ZN(\RegFile/_0280_ ) );
NAND3_X1 \RegFile/_7132_ ( .A1(\RegFile/_2606_ ), .A2(\RegFile/_2149_ ), .A3(\RegFile/_2607_ ), .ZN(\RegFile/_2878_ ) );
OAI21_X1 \RegFile/_7133_ ( .A(\RegFile/_2878_ ), .B1(\RegFile/_1891_ ), .B2(\RegFile/_2852_ ), .ZN(\RegFile/_0281_ ) );
AOI21_X1 \RegFile/_7134_ ( .A(\RegFile/_3620_ ), .B1(\RegFile/_2846_ ), .B2(\RegFile/_2848_ ), .ZN(\RegFile/_2879_ ) );
AOI21_X1 \RegFile/_7135_ ( .A(\RegFile/_2879_ ), .B1(\RegFile/_2628_ ), .B2(\RegFile/_2850_ ), .ZN(\RegFile/_0282_ ) );
NAND2_X1 \RegFile/_7136_ ( .A1(\RegFile/_2856_ ), .A2(\RegFile/_3621_ ), .ZN(\RegFile/_2880_ ) );
OAI21_X1 \RegFile/_7137_ ( .A(\RegFile/_2880_ ), .B1(\RegFile/_2646_ ), .B2(\RegFile/_2856_ ), .ZN(\RegFile/_0283_ ) );
AOI21_X1 \RegFile/_7138_ ( .A(\RegFile/_3622_ ), .B1(\RegFile/_2846_ ), .B2(\RegFile/_2848_ ), .ZN(\RegFile/_2881_ ) );
AOI21_X1 \RegFile/_7139_ ( .A(\RegFile/_2881_ ), .B1(\RegFile/_2664_ ), .B2(\RegFile/_2850_ ), .ZN(\RegFile/_0284_ ) );
AOI21_X1 \RegFile/_7140_ ( .A(\RegFile/_3623_ ), .B1(\RegFile/_2846_ ), .B2(\RegFile/_2848_ ), .ZN(\RegFile/_2882_ ) );
AOI21_X1 \RegFile/_7141_ ( .A(\RegFile/_2882_ ), .B1(\RegFile/_2685_ ), .B2(\RegFile/_2850_ ), .ZN(\RegFile/_0285_ ) );
BUF_X4 \RegFile/_7142_ ( .A(\RegFile/_2338_ ), .Z(\RegFile/_2883_ ) );
BUF_X4 \RegFile/_7143_ ( .A(\RegFile/_2847_ ), .Z(\RegFile/_2884_ ) );
AOI21_X1 \RegFile/_7144_ ( .A(\RegFile/_3625_ ), .B1(\RegFile/_2883_ ), .B2(\RegFile/_2884_ ), .ZN(\RegFile/_2885_ ) );
AOI21_X1 \RegFile/_7145_ ( .A(\RegFile/_2885_ ), .B1(\RegFile/_2705_ ), .B2(\RegFile/_2852_ ), .ZN(\RegFile/_0286_ ) );
AOI21_X1 \RegFile/_7146_ ( .A(\RegFile/_3626_ ), .B1(\RegFile/_2883_ ), .B2(\RegFile/_2884_ ), .ZN(\RegFile/_2886_ ) );
AOI21_X1 \RegFile/_7147_ ( .A(\RegFile/_2886_ ), .B1(\RegFile/_2724_ ), .B2(\RegFile/_2852_ ), .ZN(\RegFile/_0287_ ) );
BUF_X4 \RegFile/_7148_ ( .A(\RegFile/_2182_ ), .Z(\RegFile/_2887_ ) );
BUF_X4 \RegFile/_7149_ ( .A(\RegFile/_2887_ ), .Z(\RegFile/_2888_ ) );
NAND2_X1 \RegFile/_7150_ ( .A1(\RegFile/_2888_ ), .A2(\RegFile/_3634_ ), .ZN(\RegFile/_2889_ ) );
BUF_X4 \RegFile/_7151_ ( .A(\RegFile/_2887_ ), .Z(\RegFile/_2890_ ) );
OAI21_X1 \RegFile/_7152_ ( .A(\RegFile/_2889_ ), .B1(\RegFile/_2072_ ), .B2(\RegFile/_2890_ ), .ZN(\RegFile/_0288_ ) );
NAND2_X1 \RegFile/_7153_ ( .A1(\RegFile/_2888_ ), .A2(\RegFile/_3645_ ), .ZN(\RegFile/_2891_ ) );
OAI21_X1 \RegFile/_7154_ ( .A(\RegFile/_2891_ ), .B1(\RegFile/_2113_ ), .B2(\RegFile/_2890_ ), .ZN(\RegFile/_0289_ ) );
AOI21_X1 \RegFile/_7155_ ( .A(\RegFile/_3656_ ), .B1(\RegFile/_2749_ ), .B2(\RegFile/_2883_ ), .ZN(\RegFile/_2892_ ) );
BUF_X4 \RegFile/_7156_ ( .A(\RegFile/_2045_ ), .Z(\RegFile/_2893_ ) );
AOI21_X1 \RegFile/_7157_ ( .A(\RegFile/_2892_ ), .B1(\RegFile/_2142_ ), .B2(\RegFile/_2893_ ), .ZN(\RegFile/_0290_ ) );
BUF_X4 \RegFile/_7158_ ( .A(\RegFile/_2045_ ), .Z(\RegFile/_2894_ ) );
NAND3_X1 \RegFile/_7159_ ( .A1(\RegFile/_2173_ ), .A2(\RegFile/_2894_ ), .A3(\RegFile/_2174_ ), .ZN(\RegFile/_2895_ ) );
OAI21_X1 \RegFile/_7160_ ( .A(\RegFile/_2895_ ), .B1(\RegFile/_1501_ ), .B2(\RegFile/_2894_ ), .ZN(\RegFile/_0291_ ) );
OR3_X1 \RegFile/_7161_ ( .A1(\RegFile/_2196_ ), .A2(\RegFile/_2182_ ), .A3(\RegFile/_2197_ ), .ZN(\RegFile/_2896_ ) );
OAI21_X1 \RegFile/_7162_ ( .A(\RegFile/_2896_ ), .B1(\RegFile/_0902_ ), .B2(\RegFile/_2894_ ), .ZN(\RegFile/_0292_ ) );
AOI21_X1 \RegFile/_7163_ ( .A(\RegFile/_2887_ ), .B1(\RegFile/_2216_ ), .B2(\RegFile/_2217_ ), .ZN(\RegFile/_2897_ ) );
AOI21_X1 \RegFile/_7164_ ( .A(\RegFile/_2897_ ), .B1(\RegFile/_1553_ ), .B2(\RegFile/_2890_ ), .ZN(\RegFile/_0293_ ) );
BUF_X4 \RegFile/_7165_ ( .A(\RegFile/_2725_ ), .Z(\RegFile/_2898_ ) );
AOI21_X1 \RegFile/_7166_ ( .A(\RegFile/_3662_ ), .B1(\RegFile/_2898_ ), .B2(\RegFile/_2883_ ), .ZN(\RegFile/_2899_ ) );
AOI21_X1 \RegFile/_7167_ ( .A(\RegFile/_2899_ ), .B1(\RegFile/_2240_ ), .B2(\RegFile/_2893_ ), .ZN(\RegFile/_0294_ ) );
NAND3_X1 \RegFile/_7168_ ( .A1(\RegFile/_2258_ ), .A2(\RegFile/_2894_ ), .A3(\RegFile/_2259_ ), .ZN(\RegFile/_2900_ ) );
OAI21_X1 \RegFile/_7169_ ( .A(\RegFile/_2900_ ), .B1(\RegFile/_0959_ ), .B2(\RegFile/_2894_ ), .ZN(\RegFile/_0295_ ) );
AOI21_X1 \RegFile/_7170_ ( .A(\RegFile/_2887_ ), .B1(\RegFile/_2278_ ), .B2(\RegFile/_2279_ ), .ZN(\RegFile/_2901_ ) );
AOI21_X1 \RegFile/_7171_ ( .A(\RegFile/_2901_ ), .B1(\RegFile/_0977_ ), .B2(\RegFile/_2890_ ), .ZN(\RegFile/_0296_ ) );
NAND3_X1 \RegFile/_7172_ ( .A1(\RegFile/_2296_ ), .A2(\RegFile/_2045_ ), .A3(\RegFile/_2297_ ), .ZN(\RegFile/_2902_ ) );
OAI21_X1 \RegFile/_7173_ ( .A(\RegFile/_2902_ ), .B1(\RegFile/_2282_ ), .B2(\RegFile/_2894_ ), .ZN(\RegFile/_0297_ ) );
NAND3_X1 \RegFile/_7174_ ( .A1(\RegFile/_2315_ ), .A2(\RegFile/_2045_ ), .A3(\RegFile/_2316_ ), .ZN(\RegFile/_2903_ ) );
OAI21_X1 \RegFile/_7175_ ( .A(\RegFile/_2903_ ), .B1(\RegFile/_1014_ ), .B2(\RegFile/_2894_ ), .ZN(\RegFile/_0298_ ) );
OR3_X1 \RegFile/_7176_ ( .A1(\RegFile/_2333_ ), .A2(\RegFile/_2182_ ), .A3(\RegFile/_2334_ ), .ZN(\RegFile/_2904_ ) );
OAI21_X1 \RegFile/_7177_ ( .A(\RegFile/_2904_ ), .B1(\RegFile/_1661_ ), .B2(\RegFile/_2894_ ), .ZN(\RegFile/_0299_ ) );
AOI21_X1 \RegFile/_7178_ ( .A(\RegFile/_2887_ ), .B1(\RegFile/_2354_ ), .B2(\RegFile/_2355_ ), .ZN(\RegFile/_2905_ ) );
AOI21_X1 \RegFile/_7179_ ( .A(\RegFile/_2905_ ), .B1(\RegFile/_1049_ ), .B2(\RegFile/_2890_ ), .ZN(\RegFile/_0300_ ) );
AOI21_X1 \RegFile/_7180_ ( .A(\RegFile/_3638_ ), .B1(\RegFile/_2898_ ), .B2(\RegFile/_2883_ ), .ZN(\RegFile/_2906_ ) );
AOI21_X1 \RegFile/_7181_ ( .A(\RegFile/_2906_ ), .B1(\RegFile/_2379_ ), .B2(\RegFile/_2893_ ), .ZN(\RegFile/_0301_ ) );
AOI21_X1 \RegFile/_7182_ ( .A(\RegFile/_2887_ ), .B1(\RegFile/_2397_ ), .B2(\RegFile/_2398_ ), .ZN(\RegFile/_2907_ ) );
AOI21_X1 \RegFile/_7183_ ( .A(\RegFile/_2907_ ), .B1(\RegFile/_1708_ ), .B2(\RegFile/_2890_ ), .ZN(\RegFile/_0302_ ) );
BUF_X2 \RegFile/_7184_ ( .A(\RegFile/_2338_ ), .Z(\RegFile/_2908_ ) );
AOI21_X1 \RegFile/_7185_ ( .A(\RegFile/_3640_ ), .B1(\RegFile/_2898_ ), .B2(\RegFile/_2908_ ), .ZN(\RegFile/_2909_ ) );
AOI21_X1 \RegFile/_7186_ ( .A(\RegFile/_2909_ ), .B1(\RegFile/_2420_ ), .B2(\RegFile/_2893_ ), .ZN(\RegFile/_0303_ ) );
NAND2_X1 \RegFile/_7187_ ( .A1(\RegFile/_2888_ ), .A2(\RegFile/_3641_ ), .ZN(\RegFile/_2910_ ) );
OAI21_X1 \RegFile/_7188_ ( .A(\RegFile/_2910_ ), .B1(\RegFile/_2440_ ), .B2(\RegFile/_2888_ ), .ZN(\RegFile/_0304_ ) );
NAND2_X1 \RegFile/_7189_ ( .A1(\RegFile/_2888_ ), .A2(\RegFile/_3642_ ), .ZN(\RegFile/_2911_ ) );
OAI21_X1 \RegFile/_7190_ ( .A(\RegFile/_2911_ ), .B1(\RegFile/_2459_ ), .B2(\RegFile/_2888_ ), .ZN(\RegFile/_0305_ ) );
AOI21_X1 \RegFile/_7191_ ( .A(\RegFile/_3643_ ), .B1(\RegFile/_2898_ ), .B2(\RegFile/_2908_ ), .ZN(\RegFile/_2912_ ) );
AOI21_X1 \RegFile/_7192_ ( .A(\RegFile/_2912_ ), .B1(\RegFile/_2476_ ), .B2(\RegFile/_2893_ ), .ZN(\RegFile/_0306_ ) );
NAND2_X1 \RegFile/_7193_ ( .A1(\RegFile/_2888_ ), .A2(\RegFile/_3644_ ), .ZN(\RegFile/_2913_ ) );
OAI21_X1 \RegFile/_7194_ ( .A(\RegFile/_2913_ ), .B1(\RegFile/_2495_ ), .B2(\RegFile/_2888_ ), .ZN(\RegFile/_0307_ ) );
AOI21_X1 \RegFile/_7195_ ( .A(\RegFile/_3646_ ), .B1(\RegFile/_2898_ ), .B2(\RegFile/_2908_ ), .ZN(\RegFile/_2914_ ) );
AOI21_X1 \RegFile/_7196_ ( .A(\RegFile/_2914_ ), .B1(\RegFile/_2514_ ), .B2(\RegFile/_2893_ ), .ZN(\RegFile/_0308_ ) );
AOI21_X1 \RegFile/_7197_ ( .A(\RegFile/_3647_ ), .B1(\RegFile/_2898_ ), .B2(\RegFile/_2908_ ), .ZN(\RegFile/_2915_ ) );
AOI21_X1 \RegFile/_7198_ ( .A(\RegFile/_2915_ ), .B1(\RegFile/_2533_ ), .B2(\RegFile/_2893_ ), .ZN(\RegFile/_0309_ ) );
AOI21_X1 \RegFile/_7199_ ( .A(\RegFile/_3648_ ), .B1(\RegFile/_2898_ ), .B2(\RegFile/_2908_ ), .ZN(\RegFile/_2916_ ) );
AOI21_X1 \RegFile/_7200_ ( .A(\RegFile/_2916_ ), .B1(\RegFile/_2552_ ), .B2(\RegFile/_2893_ ), .ZN(\RegFile/_0310_ ) );
NAND2_X1 \RegFile/_7201_ ( .A1(\RegFile/_2888_ ), .A2(\RegFile/_3649_ ), .ZN(\RegFile/_2917_ ) );
OAI21_X1 \RegFile/_7202_ ( .A(\RegFile/_2917_ ), .B1(\RegFile/_2571_ ), .B2(\RegFile/_2888_ ), .ZN(\RegFile/_0311_ ) );
AOI21_X1 \RegFile/_7203_ ( .A(\RegFile/_3650_ ), .B1(\RegFile/_2898_ ), .B2(\RegFile/_2908_ ), .ZN(\RegFile/_2918_ ) );
AOI21_X1 \RegFile/_7204_ ( .A(\RegFile/_2918_ ), .B1(\RegFile/_2592_ ), .B2(\RegFile/_2893_ ), .ZN(\RegFile/_0312_ ) );
AOI21_X1 \RegFile/_7205_ ( .A(\RegFile/_2887_ ), .B1(\RegFile/_2606_ ), .B2(\RegFile/_2607_ ), .ZN(\RegFile/_2919_ ) );
AOI21_X1 \RegFile/_7206_ ( .A(\RegFile/_2919_ ), .B1(\RegFile/_1264_ ), .B2(\RegFile/_2890_ ), .ZN(\RegFile/_0313_ ) );
AOI21_X1 \RegFile/_7207_ ( .A(\RegFile/_2887_ ), .B1(\RegFile/_2625_ ), .B2(\RegFile/_2626_ ), .ZN(\RegFile/_2920_ ) );
AOI21_X1 \RegFile/_7208_ ( .A(\RegFile/_2920_ ), .B1(\RegFile/_1281_ ), .B2(\RegFile/_2890_ ), .ZN(\RegFile/_0314_ ) );
AOI21_X1 \RegFile/_7209_ ( .A(\RegFile/_2887_ ), .B1(\RegFile/_2643_ ), .B2(\RegFile/_2644_ ), .ZN(\RegFile/_2921_ ) );
AOI21_X1 \RegFile/_7210_ ( .A(\RegFile/_2921_ ), .B1(\RegFile/_1920_ ), .B2(\RegFile/_2890_ ), .ZN(\RegFile/_0315_ ) );
OR3_X1 \RegFile/_7211_ ( .A1(\RegFile/_2661_ ), .A2(\RegFile/_2182_ ), .A3(\RegFile/_2662_ ), .ZN(\RegFile/_2922_ ) );
OAI21_X1 \RegFile/_7212_ ( .A(\RegFile/_2922_ ), .B1(\RegFile/_1315_ ), .B2(\RegFile/_2894_ ), .ZN(\RegFile/_0316_ ) );
AOI21_X1 \RegFile/_7213_ ( .A(\RegFile/_3655_ ), .B1(\RegFile/_2898_ ), .B2(\RegFile/_2908_ ), .ZN(\RegFile/_2923_ ) );
AOI21_X1 \RegFile/_7214_ ( .A(\RegFile/_2923_ ), .B1(\RegFile/_2685_ ), .B2(\RegFile/_2893_ ), .ZN(\RegFile/_0317_ ) );
NAND3_X1 \RegFile/_7215_ ( .A1(\RegFile/_2702_ ), .A2(\RegFile/_2045_ ), .A3(\RegFile/_2703_ ), .ZN(\RegFile/_2924_ ) );
OAI21_X1 \RegFile/_7216_ ( .A(\RegFile/_2924_ ), .B1(\RegFile/_1353_ ), .B2(\RegFile/_2894_ ), .ZN(\RegFile/_0318_ ) );
AOI21_X1 \RegFile/_7217_ ( .A(\RegFile/_2887_ ), .B1(\RegFile/_2721_ ), .B2(\RegFile/_2722_ ), .ZN(\RegFile/_2925_ ) );
AOI21_X1 \RegFile/_7218_ ( .A(\RegFile/_2925_ ), .B1(\RegFile/_1378_ ), .B2(\RegFile/_2890_ ), .ZN(\RegFile/_0319_ ) );
BUF_X4 \RegFile/_7219_ ( .A(\RegFile/_2118_ ), .Z(\RegFile/_2926_ ) );
NAND2_X1 \RegFile/_7220_ ( .A1(\RegFile/_2926_ ), .A2(\RegFile/_3666_ ), .ZN(\RegFile/_2927_ ) );
BUF_X4 \RegFile/_7221_ ( .A(\RegFile/_2118_ ), .Z(\RegFile/_2928_ ) );
BUF_X4 \RegFile/_7222_ ( .A(\RegFile/_2928_ ), .Z(\RegFile/_2929_ ) );
OAI21_X1 \RegFile/_7223_ ( .A(\RegFile/_2927_ ), .B1(\RegFile/_2071_ ), .B2(\RegFile/_2929_ ), .ZN(\RegFile/_0320_ ) );
AOI21_X1 \RegFile/_7224_ ( .A(\RegFile/_2928_ ), .B1(\RegFile/_2110_ ), .B2(\RegFile/_2111_ ), .ZN(\RegFile/_2930_ ) );
BUF_X4 \RegFile/_7225_ ( .A(\RegFile/_2928_ ), .Z(\RegFile/_2931_ ) );
AOI21_X1 \RegFile/_7226_ ( .A(\RegFile/_2930_ ), .B1(\RegFile/_0817_ ), .B2(\RegFile/_2931_ ), .ZN(\RegFile/_0321_ ) );
AOI21_X1 \RegFile/_7227_ ( .A(\RegFile/_2928_ ), .B1(\RegFile/_2139_ ), .B2(\RegFile/_2140_ ), .ZN(\RegFile/_2932_ ) );
AOI21_X1 \RegFile/_7228_ ( .A(\RegFile/_2932_ ), .B1(\RegFile/_0856_ ), .B2(\RegFile/_2931_ ), .ZN(\RegFile/_0322_ ) );
NAND2_X1 \RegFile/_7229_ ( .A1(\RegFile/_2926_ ), .A2(\RegFile/_3691_ ), .ZN(\RegFile/_2933_ ) );
OAI21_X1 \RegFile/_7230_ ( .A(\RegFile/_2933_ ), .B1(\RegFile/_2175_ ), .B2(\RegFile/_2929_ ), .ZN(\RegFile/_0323_ ) );
NAND2_X1 \RegFile/_7231_ ( .A1(\RegFile/_2926_ ), .A2(\RegFile/_3692_ ), .ZN(\RegFile/_2934_ ) );
OAI21_X1 \RegFile/_7232_ ( .A(\RegFile/_2934_ ), .B1(\RegFile/_2199_ ), .B2(\RegFile/_2929_ ), .ZN(\RegFile/_0324_ ) );
NAND2_X1 \RegFile/_7233_ ( .A1(\RegFile/_2926_ ), .A2(\RegFile/_3693_ ), .ZN(\RegFile/_2935_ ) );
OAI21_X1 \RegFile/_7234_ ( .A(\RegFile/_2935_ ), .B1(\RegFile/_2218_ ), .B2(\RegFile/_2929_ ), .ZN(\RegFile/_0325_ ) );
NAND2_X1 \RegFile/_7235_ ( .A1(\RegFile/_2926_ ), .A2(\RegFile/_3694_ ), .ZN(\RegFile/_2936_ ) );
OAI21_X1 \RegFile/_7236_ ( .A(\RegFile/_2936_ ), .B1(\RegFile/_2240_ ), .B2(\RegFile/_2929_ ), .ZN(\RegFile/_0326_ ) );
NAND2_X1 \RegFile/_7237_ ( .A1(\RegFile/_2926_ ), .A2(\RegFile/_3695_ ), .ZN(\RegFile/_2937_ ) );
OAI21_X1 \RegFile/_7238_ ( .A(\RegFile/_2937_ ), .B1(\RegFile/_2260_ ), .B2(\RegFile/_2929_ ), .ZN(\RegFile/_0327_ ) );
AOI21_X1 \RegFile/_7239_ ( .A(\RegFile/_2928_ ), .B1(\RegFile/_2278_ ), .B2(\RegFile/_2279_ ), .ZN(\RegFile/_2938_ ) );
AOI21_X1 \RegFile/_7240_ ( .A(\RegFile/_2938_ ), .B1(\RegFile/_0976_ ), .B2(\RegFile/_2931_ ), .ZN(\RegFile/_0328_ ) );
AOI21_X1 \RegFile/_7241_ ( .A(\RegFile/_2928_ ), .B1(\RegFile/_2296_ ), .B2(\RegFile/_2297_ ), .ZN(\RegFile/_2939_ ) );
AOI21_X1 \RegFile/_7242_ ( .A(\RegFile/_2939_ ), .B1(\RegFile/_0996_ ), .B2(\RegFile/_2931_ ), .ZN(\RegFile/_0329_ ) );
AOI21_X1 \RegFile/_7243_ ( .A(\RegFile/_2928_ ), .B1(\RegFile/_2315_ ), .B2(\RegFile/_2316_ ), .ZN(\RegFile/_2940_ ) );
AOI21_X1 \RegFile/_7244_ ( .A(\RegFile/_2940_ ), .B1(\RegFile/_1013_ ), .B2(\RegFile/_2931_ ), .ZN(\RegFile/_0330_ ) );
NAND2_X1 \RegFile/_7245_ ( .A1(\RegFile/_2926_ ), .A2(\RegFile/_3668_ ), .ZN(\RegFile/_2941_ ) );
BUF_X4 \RegFile/_7246_ ( .A(\RegFile/_2928_ ), .Z(\RegFile/_2942_ ) );
OAI21_X1 \RegFile/_7247_ ( .A(\RegFile/_2941_ ), .B1(\RegFile/_2336_ ), .B2(\RegFile/_2942_ ), .ZN(\RegFile/_0331_ ) );
AOI21_X1 \RegFile/_7248_ ( .A(\RegFile/_2928_ ), .B1(\RegFile/_2354_ ), .B2(\RegFile/_2355_ ), .ZN(\RegFile/_2943_ ) );
AOI21_X1 \RegFile/_7249_ ( .A(\RegFile/_2943_ ), .B1(\RegFile/_1048_ ), .B2(\RegFile/_2931_ ), .ZN(\RegFile/_0332_ ) );
NAND2_X1 \RegFile/_7250_ ( .A1(\RegFile/_2926_ ), .A2(\RegFile/_3670_ ), .ZN(\RegFile/_2944_ ) );
OAI21_X1 \RegFile/_7251_ ( .A(\RegFile/_2944_ ), .B1(\RegFile/_2379_ ), .B2(\RegFile/_2942_ ), .ZN(\RegFile/_0333_ ) );
BUF_X4 \RegFile/_7252_ ( .A(\RegFile/_2118_ ), .Z(\RegFile/_2945_ ) );
NAND2_X1 \RegFile/_7253_ ( .A1(\RegFile/_2945_ ), .A2(\RegFile/_3671_ ), .ZN(\RegFile/_2946_ ) );
OAI21_X1 \RegFile/_7254_ ( .A(\RegFile/_2946_ ), .B1(\RegFile/_2399_ ), .B2(\RegFile/_2942_ ), .ZN(\RegFile/_0334_ ) );
AOI21_X1 \RegFile/_7255_ ( .A(\RegFile/_2928_ ), .B1(\RegFile/_2417_ ), .B2(\RegFile/_2418_ ), .ZN(\RegFile/_2947_ ) );
AOI21_X1 \RegFile/_7256_ ( .A(\RegFile/_2947_ ), .B1(\RegFile/_1720_ ), .B2(\RegFile/_2931_ ), .ZN(\RegFile/_0335_ ) );
AOI21_X1 \RegFile/_7257_ ( .A(\RegFile/_2118_ ), .B1(\RegFile/_2437_ ), .B2(\RegFile/_2438_ ), .ZN(\RegFile/_2948_ ) );
AOI21_X1 \RegFile/_7258_ ( .A(\RegFile/_2948_ ), .B1(\RegFile/_1735_ ), .B2(\RegFile/_2931_ ), .ZN(\RegFile/_0336_ ) );
NAND2_X1 \RegFile/_7259_ ( .A1(\RegFile/_2945_ ), .A2(\RegFile/_3674_ ), .ZN(\RegFile/_2949_ ) );
OAI21_X1 \RegFile/_7260_ ( .A(\RegFile/_2949_ ), .B1(\RegFile/_2459_ ), .B2(\RegFile/_2942_ ), .ZN(\RegFile/_0337_ ) );
AOI21_X1 \RegFile/_7261_ ( .A(\RegFile/_2118_ ), .B1(\RegFile/_2473_ ), .B2(\RegFile/_2474_ ), .ZN(\RegFile/_2950_ ) );
AOI21_X1 \RegFile/_7262_ ( .A(\RegFile/_2950_ ), .B1(\RegFile/_1155_ ), .B2(\RegFile/_2931_ ), .ZN(\RegFile/_0338_ ) );
BUF_X2 \RegFile/_7263_ ( .A(\RegFile/_2169_ ), .Z(\RegFile/_2951_ ) );
AND3_X1 \RegFile/_7264_ ( .A1(\RegFile/_2494_ ), .A2(\RegFile/_2908_ ), .A3(\RegFile/_2951_ ), .ZN(\RegFile/_2952_ ) );
AOI21_X1 \RegFile/_7265_ ( .A(\RegFile/_2952_ ), .B1(\RegFile/_1165_ ), .B2(\RegFile/_2931_ ), .ZN(\RegFile/_0339_ ) );
AND3_X4 \RegFile/_7266_ ( .A1(\RegFile/_2513_ ), .A2(\RegFile/_2908_ ), .A3(\RegFile/_2951_ ), .ZN(\RegFile/_2953_ ) );
AOI21_X1 \RegFile/_7267_ ( .A(\RegFile/_2953_ ), .B1(\RegFile/_1183_ ), .B2(\RegFile/_2929_ ), .ZN(\RegFile/_0340_ ) );
NAND2_X1 \RegFile/_7268_ ( .A1(\RegFile/_2945_ ), .A2(\RegFile/_3679_ ), .ZN(\RegFile/_2954_ ) );
OAI21_X1 \RegFile/_7269_ ( .A(\RegFile/_2954_ ), .B1(\RegFile/_2533_ ), .B2(\RegFile/_2942_ ), .ZN(\RegFile/_0341_ ) );
NAND2_X1 \RegFile/_7270_ ( .A1(\RegFile/_2945_ ), .A2(\RegFile/_3680_ ), .ZN(\RegFile/_2955_ ) );
OAI21_X1 \RegFile/_7271_ ( .A(\RegFile/_2955_ ), .B1(\RegFile/_2552_ ), .B2(\RegFile/_2942_ ), .ZN(\RegFile/_0342_ ) );
NAND2_X1 \RegFile/_7272_ ( .A1(\RegFile/_2945_ ), .A2(\RegFile/_3681_ ), .ZN(\RegFile/_2956_ ) );
OAI21_X1 \RegFile/_7273_ ( .A(\RegFile/_2956_ ), .B1(\RegFile/_2571_ ), .B2(\RegFile/_2942_ ), .ZN(\RegFile/_0343_ ) );
AOI21_X1 \RegFile/_7274_ ( .A(\RegFile/_2118_ ), .B1(\RegFile/_2589_ ), .B2(\RegFile/_2590_ ), .ZN(\RegFile/_2957_ ) );
AOI21_X1 \RegFile/_7275_ ( .A(\RegFile/_2957_ ), .B1(\RegFile/_1248_ ), .B2(\RegFile/_2929_ ), .ZN(\RegFile/_0344_ ) );
NAND2_X1 \RegFile/_7276_ ( .A1(\RegFile/_2945_ ), .A2(\RegFile/_3683_ ), .ZN(\RegFile/_2958_ ) );
OAI21_X1 \RegFile/_7277_ ( .A(\RegFile/_2958_ ), .B1(\RegFile/_2608_ ), .B2(\RegFile/_2942_ ), .ZN(\RegFile/_0345_ ) );
AOI21_X1 \RegFile/_7278_ ( .A(\RegFile/_2118_ ), .B1(\RegFile/_2625_ ), .B2(\RegFile/_2626_ ), .ZN(\RegFile/_2959_ ) );
AOI21_X1 \RegFile/_7279_ ( .A(\RegFile/_2959_ ), .B1(\RegFile/_1280_ ), .B2(\RegFile/_2929_ ), .ZN(\RegFile/_0346_ ) );
NAND2_X1 \RegFile/_7280_ ( .A1(\RegFile/_2945_ ), .A2(\RegFile/_3685_ ), .ZN(\RegFile/_2960_ ) );
OAI21_X1 \RegFile/_7281_ ( .A(\RegFile/_2960_ ), .B1(\RegFile/_2646_ ), .B2(\RegFile/_2942_ ), .ZN(\RegFile/_0347_ ) );
AND3_X4 \RegFile/_7282_ ( .A1(\RegFile/_2663_ ), .A2(\RegFile/_2908_ ), .A3(\RegFile/_2169_ ), .ZN(\RegFile/_2961_ ) );
AOI21_X1 \RegFile/_7283_ ( .A(\RegFile/_2961_ ), .B1(\RegFile/_1314_ ), .B2(\RegFile/_2929_ ), .ZN(\RegFile/_0348_ ) );
NAND2_X1 \RegFile/_7284_ ( .A1(\RegFile/_2945_ ), .A2(\RegFile/_3687_ ), .ZN(\RegFile/_2962_ ) );
OAI21_X1 \RegFile/_7285_ ( .A(\RegFile/_2962_ ), .B1(\RegFile/_2684_ ), .B2(\RegFile/_2942_ ), .ZN(\RegFile/_0349_ ) );
NAND2_X1 \RegFile/_7286_ ( .A1(\RegFile/_2945_ ), .A2(\RegFile/_3689_ ), .ZN(\RegFile/_2963_ ) );
OAI21_X1 \RegFile/_7287_ ( .A(\RegFile/_2963_ ), .B1(\RegFile/_2705_ ), .B2(\RegFile/_2926_ ), .ZN(\RegFile/_0350_ ) );
NAND2_X1 \RegFile/_7288_ ( .A1(\RegFile/_2945_ ), .A2(\RegFile/_3690_ ), .ZN(\RegFile/_2964_ ) );
OAI21_X1 \RegFile/_7289_ ( .A(\RegFile/_2964_ ), .B1(\RegFile/_2723_ ), .B2(\RegFile/_2926_ ), .ZN(\RegFile/_0351_ ) );
BUF_X4 \RegFile/_7290_ ( .A(\RegFile/_2116_ ), .Z(\RegFile/_2965_ ) );
BUF_X4 \RegFile/_7291_ ( .A(\RegFile/_2965_ ), .Z(\RegFile/_2966_ ) );
NAND2_X1 \RegFile/_7292_ ( .A1(\RegFile/_2966_ ), .A2(\RegFile/_3698_ ), .ZN(\RegFile/_2967_ ) );
BUF_X4 \RegFile/_7293_ ( .A(\RegFile/_2965_ ), .Z(\RegFile/_2968_ ) );
OAI21_X1 \RegFile/_7294_ ( .A(\RegFile/_2967_ ), .B1(\RegFile/_2071_ ), .B2(\RegFile/_2968_ ), .ZN(\RegFile/_0352_ ) );
BUF_X4 \RegFile/_7295_ ( .A(\RegFile/_2152_ ), .Z(\RegFile/_2969_ ) );
NAND3_X1 \RegFile/_7296_ ( .A1(\RegFile/_2110_ ), .A2(\RegFile/_2969_ ), .A3(\RegFile/_2111_ ), .ZN(\RegFile/_2970_ ) );
BUF_X4 \RegFile/_7297_ ( .A(\RegFile/_2152_ ), .Z(\RegFile/_2971_ ) );
BUF_X4 \RegFile/_7298_ ( .A(\RegFile/_2971_ ), .Z(\RegFile/_2972_ ) );
OAI21_X1 \RegFile/_7299_ ( .A(\RegFile/_2970_ ), .B1(\RegFile/_0849_ ), .B2(\RegFile/_2972_ ), .ZN(\RegFile/_0353_ ) );
NAND3_X1 \RegFile/_7300_ ( .A1(\RegFile/_2139_ ), .A2(\RegFile/_2971_ ), .A3(\RegFile/_2140_ ), .ZN(\RegFile/_2973_ ) );
OAI21_X1 \RegFile/_7301_ ( .A(\RegFile/_2973_ ), .B1(\RegFile/_0859_ ), .B2(\RegFile/_2972_ ), .ZN(\RegFile/_0354_ ) );
NAND3_X1 \RegFile/_7302_ ( .A1(\RegFile/_2173_ ), .A2(\RegFile/_2971_ ), .A3(\RegFile/_2174_ ), .ZN(\RegFile/_2974_ ) );
OAI21_X1 \RegFile/_7303_ ( .A(\RegFile/_2974_ ), .B1(\RegFile/_1515_ ), .B2(\RegFile/_2972_ ), .ZN(\RegFile/_0355_ ) );
AND2_X1 \RegFile/_7304_ ( .A1(\RegFile/_2198_ ), .A2(\RegFile/_2152_ ), .ZN(\RegFile/_2975_ ) );
AOI21_X1 \RegFile/_7305_ ( .A(\RegFile/_2975_ ), .B1(\RegFile/_0905_ ), .B2(\RegFile/_2968_ ), .ZN(\RegFile/_0356_ ) );
NAND3_X1 \RegFile/_7306_ ( .A1(\RegFile/_2216_ ), .A2(\RegFile/_2971_ ), .A3(\RegFile/_2217_ ), .ZN(\RegFile/_2976_ ) );
OAI21_X1 \RegFile/_7307_ ( .A(\RegFile/_2976_ ), .B1(\RegFile/_1549_ ), .B2(\RegFile/_2972_ ), .ZN(\RegFile/_0357_ ) );
AOI21_X1 \RegFile/_7308_ ( .A(\RegFile/_2965_ ), .B1(\RegFile/_2235_ ), .B2(\RegFile/_2238_ ), .ZN(\RegFile/_2977_ ) );
AOI21_X1 \RegFile/_7309_ ( .A(\RegFile/_2977_ ), .B1(\RegFile/_1574_ ), .B2(\RegFile/_2968_ ), .ZN(\RegFile/_0358_ ) );
AOI21_X1 \RegFile/_7310_ ( .A(\RegFile/_3727_ ), .B1(\RegFile/_2883_ ), .B2(\RegFile/_2839_ ), .ZN(\RegFile/_2978_ ) );
AOI21_X1 \RegFile/_7311_ ( .A(\RegFile/_2978_ ), .B1(\RegFile/_2261_ ), .B2(\RegFile/_2972_ ), .ZN(\RegFile/_0359_ ) );
AOI21_X1 \RegFile/_7312_ ( .A(\RegFile/_3728_ ), .B1(\RegFile/_2883_ ), .B2(\RegFile/_2839_ ), .ZN(\RegFile/_2979_ ) );
AOI21_X1 \RegFile/_7313_ ( .A(\RegFile/_2979_ ), .B1(\RegFile/_2782_ ), .B2(\RegFile/_2972_ ), .ZN(\RegFile/_0360_ ) );
AOI21_X1 \RegFile/_7314_ ( .A(\RegFile/_2965_ ), .B1(\RegFile/_2296_ ), .B2(\RegFile/_2297_ ), .ZN(\RegFile/_2980_ ) );
AOI21_X1 \RegFile/_7315_ ( .A(\RegFile/_2980_ ), .B1(\RegFile/_1009_ ), .B2(\RegFile/_2968_ ), .ZN(\RegFile/_0361_ ) );
NAND2_X1 \RegFile/_7316_ ( .A1(\RegFile/_2966_ ), .A2(\RegFile/_3699_ ), .ZN(\RegFile/_2981_ ) );
OAI21_X1 \RegFile/_7317_ ( .A(\RegFile/_2981_ ), .B1(\RegFile/_2317_ ), .B2(\RegFile/_2968_ ), .ZN(\RegFile/_0362_ ) );
AND2_X1 \RegFile/_7318_ ( .A1(\RegFile/_2335_ ), .A2(\RegFile/_2152_ ), .ZN(\RegFile/_2982_ ) );
AOI21_X1 \RegFile/_7319_ ( .A(\RegFile/_2982_ ), .B1(\RegFile/_1657_ ), .B2(\RegFile/_2968_ ), .ZN(\RegFile/_0363_ ) );
NAND3_X1 \RegFile/_7320_ ( .A1(\RegFile/_2354_ ), .A2(\RegFile/_2971_ ), .A3(\RegFile/_2355_ ), .ZN(\RegFile/_2983_ ) );
OAI21_X1 \RegFile/_7321_ ( .A(\RegFile/_2983_ ), .B1(\RegFile/_1052_ ), .B2(\RegFile/_2972_ ), .ZN(\RegFile/_0364_ ) );
AOI21_X1 \RegFile/_7322_ ( .A(\RegFile/_3702_ ), .B1(\RegFile/_2883_ ), .B2(\RegFile/_2839_ ), .ZN(\RegFile/_2984_ ) );
AOI21_X1 \RegFile/_7323_ ( .A(\RegFile/_2984_ ), .B1(\RegFile/_2379_ ), .B2(\RegFile/_2972_ ), .ZN(\RegFile/_0365_ ) );
NAND3_X1 \RegFile/_7324_ ( .A1(\RegFile/_2397_ ), .A2(\RegFile/_2971_ ), .A3(\RegFile/_2398_ ), .ZN(\RegFile/_2985_ ) );
OAI21_X1 \RegFile/_7325_ ( .A(\RegFile/_2985_ ), .B1(\RegFile/_1705_ ), .B2(\RegFile/_2969_ ), .ZN(\RegFile/_0366_ ) );
NAND2_X1 \RegFile/_7326_ ( .A1(\RegFile/_2966_ ), .A2(\RegFile/_3704_ ), .ZN(\RegFile/_2986_ ) );
OAI21_X1 \RegFile/_7327_ ( .A(\RegFile/_2986_ ), .B1(\RegFile/_2420_ ), .B2(\RegFile/_2968_ ), .ZN(\RegFile/_0367_ ) );
NAND2_X1 \RegFile/_7328_ ( .A1(\RegFile/_2966_ ), .A2(\RegFile/_3705_ ), .ZN(\RegFile/_2987_ ) );
OAI21_X1 \RegFile/_7329_ ( .A(\RegFile/_2987_ ), .B1(\RegFile/_2440_ ), .B2(\RegFile/_2968_ ), .ZN(\RegFile/_0368_ ) );
OR3_X1 \RegFile/_7330_ ( .A1(\RegFile/_2456_ ), .A2(\RegFile/_2965_ ), .A3(\RegFile/_2457_ ), .ZN(\RegFile/_2988_ ) );
OAI21_X1 \RegFile/_7331_ ( .A(\RegFile/_2988_ ), .B1(\RegFile/_1141_ ), .B2(\RegFile/_2969_ ), .ZN(\RegFile/_0369_ ) );
AOI21_X1 \RegFile/_7332_ ( .A(\RegFile/_2965_ ), .B1(\RegFile/_2473_ ), .B2(\RegFile/_2474_ ), .ZN(\RegFile/_2989_ ) );
AOI21_X1 \RegFile/_7333_ ( .A(\RegFile/_2989_ ), .B1(\RegFile/_1158_ ), .B2(\RegFile/_2968_ ), .ZN(\RegFile/_0370_ ) );
OR3_X1 \RegFile/_7334_ ( .A1(\RegFile/_2492_ ), .A2(\RegFile/_2965_ ), .A3(\RegFile/_2493_ ), .ZN(\RegFile/_2990_ ) );
OAI21_X1 \RegFile/_7335_ ( .A(\RegFile/_2990_ ), .B1(\RegFile/_1178_ ), .B2(\RegFile/_2969_ ), .ZN(\RegFile/_0371_ ) );
OR3_X1 \RegFile/_7336_ ( .A1(\RegFile/_2511_ ), .A2(\RegFile/_2965_ ), .A3(\RegFile/_2512_ ), .ZN(\RegFile/_2991_ ) );
OAI21_X1 \RegFile/_7337_ ( .A(\RegFile/_2991_ ), .B1(\RegFile/_1187_ ), .B2(\RegFile/_2969_ ), .ZN(\RegFile/_0372_ ) );
NAND3_X1 \RegFile/_7338_ ( .A1(\RegFile/_2530_ ), .A2(\RegFile/_2971_ ), .A3(\RegFile/_2531_ ), .ZN(\RegFile/_2992_ ) );
OAI21_X1 \RegFile/_7339_ ( .A(\RegFile/_2992_ ), .B1(\RegFile/_1819_ ), .B2(\RegFile/_2969_ ), .ZN(\RegFile/_0373_ ) );
AOI21_X1 \RegFile/_7340_ ( .A(\RegFile/_2965_ ), .B1(\RegFile/_2549_ ), .B2(\RegFile/_2550_ ), .ZN(\RegFile/_2993_ ) );
AOI21_X1 \RegFile/_7341_ ( .A(\RegFile/_2993_ ), .B1(\RegFile/_1838_ ), .B2(\RegFile/_2968_ ), .ZN(\RegFile/_0374_ ) );
NAND3_X1 \RegFile/_7342_ ( .A1(\RegFile/_2568_ ), .A2(\RegFile/_2971_ ), .A3(\RegFile/_2569_ ), .ZN(\RegFile/_2994_ ) );
OAI21_X1 \RegFile/_7343_ ( .A(\RegFile/_2994_ ), .B1(\RegFile/_1858_ ), .B2(\RegFile/_2969_ ), .ZN(\RegFile/_0375_ ) );
NAND2_X1 \RegFile/_7344_ ( .A1(\RegFile/_2966_ ), .A2(\RegFile/_3714_ ), .ZN(\RegFile/_2995_ ) );
OAI21_X1 \RegFile/_7345_ ( .A(\RegFile/_2995_ ), .B1(\RegFile/_2592_ ), .B2(\RegFile/_2966_ ), .ZN(\RegFile/_0376_ ) );
NAND3_X1 \RegFile/_7346_ ( .A1(\RegFile/_2606_ ), .A2(\RegFile/_2971_ ), .A3(\RegFile/_2607_ ), .ZN(\RegFile/_2996_ ) );
OAI21_X1 \RegFile/_7347_ ( .A(\RegFile/_2996_ ), .B1(\RegFile/_1275_ ), .B2(\RegFile/_2969_ ), .ZN(\RegFile/_0377_ ) );
NAND2_X1 \RegFile/_7348_ ( .A1(\RegFile/_2966_ ), .A2(\RegFile/_3716_ ), .ZN(\RegFile/_2997_ ) );
OAI21_X1 \RegFile/_7349_ ( .A(\RegFile/_2997_ ), .B1(\RegFile/_2627_ ), .B2(\RegFile/_2966_ ), .ZN(\RegFile/_0378_ ) );
NAND3_X1 \RegFile/_7350_ ( .A1(\RegFile/_2643_ ), .A2(\RegFile/_2971_ ), .A3(\RegFile/_2644_ ), .ZN(\RegFile/_2998_ ) );
OAI21_X1 \RegFile/_7351_ ( .A(\RegFile/_2998_ ), .B1(\RegFile/_1916_ ), .B2(\RegFile/_2969_ ), .ZN(\RegFile/_0379_ ) );
OR3_X1 \RegFile/_7352_ ( .A1(\RegFile/_2661_ ), .A2(\RegFile/_2965_ ), .A3(\RegFile/_2662_ ), .ZN(\RegFile/_2999_ ) );
OAI21_X1 \RegFile/_7353_ ( .A(\RegFile/_2999_ ), .B1(\RegFile/_1318_ ), .B2(\RegFile/_2969_ ), .ZN(\RegFile/_0380_ ) );
AOI21_X1 \RegFile/_7354_ ( .A(\RegFile/_3719_ ), .B1(\RegFile/_2883_ ), .B2(\RegFile/_2839_ ), .ZN(\RegFile/_3000_ ) );
AOI21_X1 \RegFile/_7355_ ( .A(\RegFile/_3000_ ), .B1(\RegFile/_2685_ ), .B2(\RegFile/_2972_ ), .ZN(\RegFile/_0381_ ) );
AOI21_X1 \RegFile/_7356_ ( .A(\RegFile/_3721_ ), .B1(\RegFile/_2883_ ), .B2(\RegFile/_2839_ ), .ZN(\RegFile/_3001_ ) );
AOI21_X1 \RegFile/_7357_ ( .A(\RegFile/_3001_ ), .B1(\RegFile/_2705_ ), .B2(\RegFile/_2972_ ), .ZN(\RegFile/_0382_ ) );
NAND2_X1 \RegFile/_7358_ ( .A1(\RegFile/_2966_ ), .A2(\RegFile/_3722_ ), .ZN(\RegFile/_3002_ ) );
OAI21_X1 \RegFile/_7359_ ( .A(\RegFile/_3002_ ), .B1(\RegFile/_2723_ ), .B2(\RegFile/_2966_ ), .ZN(\RegFile/_0383_ ) );
INV_X1 \RegFile/_7360_ ( .A(\RegFile/_2005_ ), .ZN(\RegFile/_3003_ ) );
BUF_X4 \RegFile/_7361_ ( .A(\RegFile/_3003_ ), .Z(\RegFile/_3004_ ) );
NAND2_X1 \RegFile/_7362_ ( .A1(\RegFile/_3004_ ), .A2(\RegFile/_3730_ ), .ZN(\RegFile/_3005_ ) );
OAI21_X1 \RegFile/_7363_ ( .A(\RegFile/_3005_ ), .B1(\RegFile/_2071_ ), .B2(\RegFile/_3004_ ), .ZN(\RegFile/_0384_ ) );
BUF_X4 \RegFile/_7364_ ( .A(\RegFile/_2160_ ), .Z(\RegFile/_3006_ ) );
BUF_X4 \RegFile/_7365_ ( .A(\RegFile/_3006_ ), .Z(\RegFile/_3007_ ) );
AOI21_X1 \RegFile/_7366_ ( .A(\RegFile/_3741_ ), .B1(\RegFile/_3007_ ), .B2(\RegFile/_2884_ ), .ZN(\RegFile/_3008_ ) );
BUF_X4 \RegFile/_7367_ ( .A(\RegFile/_2005_ ), .Z(\RegFile/_3009_ ) );
AOI21_X1 \RegFile/_7368_ ( .A(\RegFile/_3008_ ), .B1(\RegFile/_2113_ ), .B2(\RegFile/_3009_ ), .ZN(\RegFile/_0385_ ) );
AOI21_X1 \RegFile/_7369_ ( .A(\RegFile/_3752_ ), .B1(\RegFile/_3007_ ), .B2(\RegFile/_2884_ ), .ZN(\RegFile/_3010_ ) );
AOI21_X1 \RegFile/_7370_ ( .A(\RegFile/_3010_ ), .B1(\RegFile/_2142_ ), .B2(\RegFile/_3009_ ), .ZN(\RegFile/_0386_ ) );
NAND2_X1 \RegFile/_7371_ ( .A1(\RegFile/_3004_ ), .A2(\RegFile/_3755_ ), .ZN(\RegFile/_3011_ ) );
OAI21_X1 \RegFile/_7372_ ( .A(\RegFile/_3011_ ), .B1(\RegFile/_2175_ ), .B2(\RegFile/_3004_ ), .ZN(\RegFile/_0387_ ) );
NAND2_X1 \RegFile/_7373_ ( .A1(\RegFile/_3004_ ), .A2(\RegFile/_3756_ ), .ZN(\RegFile/_3012_ ) );
OAI21_X1 \RegFile/_7374_ ( .A(\RegFile/_3012_ ), .B1(\RegFile/_2199_ ), .B2(\RegFile/_3004_ ), .ZN(\RegFile/_0388_ ) );
AOI21_X1 \RegFile/_7375_ ( .A(\RegFile/_3757_ ), .B1(\RegFile/_3007_ ), .B2(\RegFile/_2884_ ), .ZN(\RegFile/_3013_ ) );
AOI21_X1 \RegFile/_7376_ ( .A(\RegFile/_3013_ ), .B1(\RegFile/_2218_ ), .B2(\RegFile/_3009_ ), .ZN(\RegFile/_0389_ ) );
AOI21_X1 \RegFile/_7377_ ( .A(\RegFile/_3758_ ), .B1(\RegFile/_3007_ ), .B2(\RegFile/_2884_ ), .ZN(\RegFile/_3014_ ) );
AOI21_X1 \RegFile/_7378_ ( .A(\RegFile/_3014_ ), .B1(\RegFile/_2240_ ), .B2(\RegFile/_3009_ ), .ZN(\RegFile/_0390_ ) );
AOI21_X1 \RegFile/_7379_ ( .A(\RegFile/_3759_ ), .B1(\RegFile/_3007_ ), .B2(\RegFile/_2884_ ), .ZN(\RegFile/_3015_ ) );
AOI21_X1 \RegFile/_7380_ ( .A(\RegFile/_3015_ ), .B1(\RegFile/_2261_ ), .B2(\RegFile/_3009_ ), .ZN(\RegFile/_0391_ ) );
AOI21_X1 \RegFile/_7381_ ( .A(\RegFile/_3760_ ), .B1(\RegFile/_3007_ ), .B2(\RegFile/_2884_ ), .ZN(\RegFile/_3016_ ) );
AOI21_X1 \RegFile/_7382_ ( .A(\RegFile/_3016_ ), .B1(\RegFile/_2782_ ), .B2(\RegFile/_3009_ ), .ZN(\RegFile/_0392_ ) );
AOI21_X1 \RegFile/_7383_ ( .A(\RegFile/_3761_ ), .B1(\RegFile/_3007_ ), .B2(\RegFile/_2884_ ), .ZN(\RegFile/_3017_ ) );
AOI21_X1 \RegFile/_7384_ ( .A(\RegFile/_3017_ ), .B1(\RegFile/_2299_ ), .B2(\RegFile/_3009_ ), .ZN(\RegFile/_0393_ ) );
AOI21_X1 \RegFile/_7385_ ( .A(\RegFile/_3731_ ), .B1(\RegFile/_3007_ ), .B2(\RegFile/_2884_ ), .ZN(\RegFile/_3018_ ) );
AOI21_X1 \RegFile/_7386_ ( .A(\RegFile/_3018_ ), .B1(\RegFile/_2318_ ), .B2(\RegFile/_3009_ ), .ZN(\RegFile/_0394_ ) );
BUF_X4 \RegFile/_7387_ ( .A(\RegFile/_2035_ ), .Z(\RegFile/_3019_ ) );
AOI21_X1 \RegFile/_7388_ ( .A(\RegFile/_3732_ ), .B1(\RegFile/_3007_ ), .B2(\RegFile/_3019_ ), .ZN(\RegFile/_3020_ ) );
AOI21_X1 \RegFile/_7389_ ( .A(\RegFile/_3020_ ), .B1(\RegFile/_2336_ ), .B2(\RegFile/_3009_ ), .ZN(\RegFile/_0395_ ) );
AOI21_X1 \RegFile/_7390_ ( .A(\RegFile/_3733_ ), .B1(\RegFile/_3007_ ), .B2(\RegFile/_3019_ ), .ZN(\RegFile/_3021_ ) );
AOI21_X1 \RegFile/_7391_ ( .A(\RegFile/_3021_ ), .B1(\RegFile/_2356_ ), .B2(\RegFile/_3009_ ), .ZN(\RegFile/_0396_ ) );
BUF_X4 \RegFile/_7392_ ( .A(\RegFile/_3006_ ), .Z(\RegFile/_3022_ ) );
AOI21_X1 \RegFile/_7393_ ( .A(\RegFile/_3734_ ), .B1(\RegFile/_3022_ ), .B2(\RegFile/_3019_ ), .ZN(\RegFile/_3023_ ) );
BUF_X4 \RegFile/_7394_ ( .A(\RegFile/_2005_ ), .Z(\RegFile/_3024_ ) );
AOI21_X1 \RegFile/_7395_ ( .A(\RegFile/_3023_ ), .B1(\RegFile/_2379_ ), .B2(\RegFile/_3024_ ), .ZN(\RegFile/_0397_ ) );
AOI21_X1 \RegFile/_7396_ ( .A(\RegFile/_3735_ ), .B1(\RegFile/_3022_ ), .B2(\RegFile/_3019_ ), .ZN(\RegFile/_3025_ ) );
AOI21_X1 \RegFile/_7397_ ( .A(\RegFile/_3025_ ), .B1(\RegFile/_2399_ ), .B2(\RegFile/_3024_ ), .ZN(\RegFile/_0398_ ) );
AOI21_X1 \RegFile/_7398_ ( .A(\RegFile/_3736_ ), .B1(\RegFile/_3022_ ), .B2(\RegFile/_3019_ ), .ZN(\RegFile/_3026_ ) );
AOI21_X1 \RegFile/_7399_ ( .A(\RegFile/_3026_ ), .B1(\RegFile/_2420_ ), .B2(\RegFile/_3024_ ), .ZN(\RegFile/_0399_ ) );
AOI21_X1 \RegFile/_7400_ ( .A(\RegFile/_3737_ ), .B1(\RegFile/_3022_ ), .B2(\RegFile/_3019_ ), .ZN(\RegFile/_3027_ ) );
AOI21_X1 \RegFile/_7401_ ( .A(\RegFile/_3027_ ), .B1(\RegFile/_2440_ ), .B2(\RegFile/_3024_ ), .ZN(\RegFile/_0400_ ) );
AOI21_X1 \RegFile/_7402_ ( .A(\RegFile/_3738_ ), .B1(\RegFile/_3022_ ), .B2(\RegFile/_3019_ ), .ZN(\RegFile/_3028_ ) );
AOI21_X1 \RegFile/_7403_ ( .A(\RegFile/_3028_ ), .B1(\RegFile/_2459_ ), .B2(\RegFile/_3024_ ), .ZN(\RegFile/_0401_ ) );
AOI21_X1 \RegFile/_7404_ ( .A(\RegFile/_3739_ ), .B1(\RegFile/_3022_ ), .B2(\RegFile/_3019_ ), .ZN(\RegFile/_3029_ ) );
AOI21_X1 \RegFile/_7405_ ( .A(\RegFile/_3029_ ), .B1(\RegFile/_2476_ ), .B2(\RegFile/_3024_ ), .ZN(\RegFile/_0402_ ) );
AOI21_X1 \RegFile/_7406_ ( .A(\RegFile/_3740_ ), .B1(\RegFile/_3022_ ), .B2(\RegFile/_3019_ ), .ZN(\RegFile/_3030_ ) );
AOI21_X1 \RegFile/_7407_ ( .A(\RegFile/_3030_ ), .B1(\RegFile/_2495_ ), .B2(\RegFile/_3024_ ), .ZN(\RegFile/_0403_ ) );
NAND2_X1 \RegFile/_7408_ ( .A1(\RegFile/_3003_ ), .A2(\RegFile/_3742_ ), .ZN(\RegFile/_3031_ ) );
OAI21_X1 \RegFile/_7409_ ( .A(\RegFile/_3031_ ), .B1(\RegFile/_2514_ ), .B2(\RegFile/_3004_ ), .ZN(\RegFile/_0404_ ) );
NAND2_X1 \RegFile/_7410_ ( .A1(\RegFile/_3003_ ), .A2(\RegFile/_3743_ ), .ZN(\RegFile/_3032_ ) );
OAI21_X1 \RegFile/_7411_ ( .A(\RegFile/_3032_ ), .B1(\RegFile/_2533_ ), .B2(\RegFile/_3004_ ), .ZN(\RegFile/_0405_ ) );
NAND2_X1 \RegFile/_7412_ ( .A1(\RegFile/_3003_ ), .A2(\RegFile/_3744_ ), .ZN(\RegFile/_3033_ ) );
OAI21_X1 \RegFile/_7413_ ( .A(\RegFile/_3033_ ), .B1(\RegFile/_2552_ ), .B2(\RegFile/_3004_ ), .ZN(\RegFile/_0406_ ) );
AOI21_X1 \RegFile/_7414_ ( .A(\RegFile/_3745_ ), .B1(\RegFile/_3022_ ), .B2(\RegFile/_3019_ ), .ZN(\RegFile/_3034_ ) );
AOI21_X1 \RegFile/_7415_ ( .A(\RegFile/_3034_ ), .B1(\RegFile/_2571_ ), .B2(\RegFile/_3024_ ), .ZN(\RegFile/_0407_ ) );
BUF_X4 \RegFile/_7416_ ( .A(\RegFile/_2035_ ), .Z(\RegFile/_3035_ ) );
AOI21_X1 \RegFile/_7417_ ( .A(\RegFile/_3746_ ), .B1(\RegFile/_3022_ ), .B2(\RegFile/_3035_ ), .ZN(\RegFile/_3036_ ) );
AOI21_X1 \RegFile/_7418_ ( .A(\RegFile/_3036_ ), .B1(\RegFile/_2592_ ), .B2(\RegFile/_3024_ ), .ZN(\RegFile/_0408_ ) );
AOI21_X1 \RegFile/_7419_ ( .A(\RegFile/_3747_ ), .B1(\RegFile/_3022_ ), .B2(\RegFile/_3035_ ), .ZN(\RegFile/_3037_ ) );
AOI21_X1 \RegFile/_7420_ ( .A(\RegFile/_3037_ ), .B1(\RegFile/_2608_ ), .B2(\RegFile/_3024_ ), .ZN(\RegFile/_0409_ ) );
BUF_X4 \RegFile/_7421_ ( .A(\RegFile/_3006_ ), .Z(\RegFile/_3038_ ) );
AOI21_X1 \RegFile/_7422_ ( .A(\RegFile/_3748_ ), .B1(\RegFile/_3038_ ), .B2(\RegFile/_3035_ ), .ZN(\RegFile/_3039_ ) );
AOI21_X1 \RegFile/_7423_ ( .A(\RegFile/_3039_ ), .B1(\RegFile/_2628_ ), .B2(\RegFile/_2005_ ), .ZN(\RegFile/_0410_ ) );
AOI21_X1 \RegFile/_7424_ ( .A(\RegFile/_3749_ ), .B1(\RegFile/_3038_ ), .B2(\RegFile/_3035_ ), .ZN(\RegFile/_3040_ ) );
AOI21_X1 \RegFile/_7425_ ( .A(\RegFile/_3040_ ), .B1(\RegFile/_2646_ ), .B2(\RegFile/_2005_ ), .ZN(\RegFile/_0411_ ) );
NAND2_X1 \RegFile/_7426_ ( .A1(\RegFile/_3003_ ), .A2(\RegFile/_3750_ ), .ZN(\RegFile/_3041_ ) );
OAI21_X1 \RegFile/_7427_ ( .A(\RegFile/_3041_ ), .B1(\RegFile/_2664_ ), .B2(\RegFile/_3004_ ), .ZN(\RegFile/_0412_ ) );
AOI21_X1 \RegFile/_7428_ ( .A(\RegFile/_3751_ ), .B1(\RegFile/_3038_ ), .B2(\RegFile/_3035_ ), .ZN(\RegFile/_3042_ ) );
AOI21_X1 \RegFile/_7429_ ( .A(\RegFile/_3042_ ), .B1(\RegFile/_2685_ ), .B2(\RegFile/_2005_ ), .ZN(\RegFile/_0413_ ) );
AOI21_X1 \RegFile/_7430_ ( .A(\RegFile/_3753_ ), .B1(\RegFile/_3038_ ), .B2(\RegFile/_3035_ ), .ZN(\RegFile/_3043_ ) );
AOI21_X1 \RegFile/_7431_ ( .A(\RegFile/_3043_ ), .B1(\RegFile/_2705_ ), .B2(\RegFile/_2005_ ), .ZN(\RegFile/_0414_ ) );
AOI21_X1 \RegFile/_7432_ ( .A(\RegFile/_3754_ ), .B1(\RegFile/_3038_ ), .B2(\RegFile/_3035_ ), .ZN(\RegFile/_3044_ ) );
AOI21_X1 \RegFile/_7433_ ( .A(\RegFile/_3044_ ), .B1(\RegFile/_2724_ ), .B2(\RegFile/_2005_ ), .ZN(\RegFile/_0415_ ) );
BUF_X4 \RegFile/_7434_ ( .A(\RegFile/_2161_ ), .Z(\RegFile/_3045_ ) );
AOI21_X1 \RegFile/_7435_ ( .A(\RegFile/_3762_ ), .B1(\RegFile/_3038_ ), .B2(\RegFile/_3045_ ), .ZN(\RegFile/_3046_ ) );
BUF_X4 \RegFile/_7436_ ( .A(\RegFile/_2014_ ), .Z(\RegFile/_3047_ ) );
AOI21_X1 \RegFile/_7437_ ( .A(\RegFile/_3046_ ), .B1(\RegFile/_2072_ ), .B2(\RegFile/_3047_ ), .ZN(\RegFile/_0416_ ) );
AOI21_X1 \RegFile/_7438_ ( .A(\RegFile/_3773_ ), .B1(\RegFile/_3038_ ), .B2(\RegFile/_3045_ ), .ZN(\RegFile/_3048_ ) );
AOI21_X1 \RegFile/_7439_ ( .A(\RegFile/_3048_ ), .B1(\RegFile/_2113_ ), .B2(\RegFile/_3047_ ), .ZN(\RegFile/_0417_ ) );
AOI21_X1 \RegFile/_7440_ ( .A(\RegFile/_3784_ ), .B1(\RegFile/_3038_ ), .B2(\RegFile/_3045_ ), .ZN(\RegFile/_3049_ ) );
AOI21_X1 \RegFile/_7441_ ( .A(\RegFile/_3049_ ), .B1(\RegFile/_2142_ ), .B2(\RegFile/_3047_ ), .ZN(\RegFile/_0418_ ) );
AOI21_X1 \RegFile/_7442_ ( .A(\RegFile/_3787_ ), .B1(\RegFile/_3038_ ), .B2(\RegFile/_3045_ ), .ZN(\RegFile/_3050_ ) );
AOI21_X1 \RegFile/_7443_ ( .A(\RegFile/_3050_ ), .B1(\RegFile/_2175_ ), .B2(\RegFile/_3047_ ), .ZN(\RegFile/_0419_ ) );
INV_X1 \RegFile/_7444_ ( .A(\RegFile/_2014_ ), .ZN(\RegFile/_3051_ ) );
BUF_X4 \RegFile/_7445_ ( .A(\RegFile/_3051_ ), .Z(\RegFile/_3052_ ) );
NAND2_X1 \RegFile/_7446_ ( .A1(\RegFile/_3052_ ), .A2(\RegFile/_3788_ ), .ZN(\RegFile/_3053_ ) );
BUF_X4 \RegFile/_7447_ ( .A(\RegFile/_3051_ ), .Z(\RegFile/_3054_ ) );
OAI21_X1 \RegFile/_7448_ ( .A(\RegFile/_3053_ ), .B1(\RegFile/_2199_ ), .B2(\RegFile/_3054_ ), .ZN(\RegFile/_0420_ ) );
NAND2_X1 \RegFile/_7449_ ( .A1(\RegFile/_3052_ ), .A2(\RegFile/_3789_ ), .ZN(\RegFile/_3055_ ) );
OAI21_X1 \RegFile/_7450_ ( .A(\RegFile/_3055_ ), .B1(\RegFile/_2218_ ), .B2(\RegFile/_3054_ ), .ZN(\RegFile/_0421_ ) );
AOI21_X1 \RegFile/_7451_ ( .A(\RegFile/_3790_ ), .B1(\RegFile/_3038_ ), .B2(\RegFile/_3045_ ), .ZN(\RegFile/_3056_ ) );
AOI21_X1 \RegFile/_7452_ ( .A(\RegFile/_3056_ ), .B1(\RegFile/_2240_ ), .B2(\RegFile/_3047_ ), .ZN(\RegFile/_0422_ ) );
BUF_X4 \RegFile/_7453_ ( .A(\RegFile/_3006_ ), .Z(\RegFile/_3057_ ) );
BUF_X4 \RegFile/_7454_ ( .A(\RegFile/_2161_ ), .Z(\RegFile/_3058_ ) );
AOI21_X1 \RegFile/_7455_ ( .A(\RegFile/_3791_ ), .B1(\RegFile/_3057_ ), .B2(\RegFile/_3058_ ), .ZN(\RegFile/_3059_ ) );
AOI21_X1 \RegFile/_7456_ ( .A(\RegFile/_3059_ ), .B1(\RegFile/_2261_ ), .B2(\RegFile/_3047_ ), .ZN(\RegFile/_0423_ ) );
AOI21_X1 \RegFile/_7457_ ( .A(\RegFile/_3792_ ), .B1(\RegFile/_3057_ ), .B2(\RegFile/_3058_ ), .ZN(\RegFile/_3060_ ) );
AOI21_X1 \RegFile/_7458_ ( .A(\RegFile/_3060_ ), .B1(\RegFile/_2782_ ), .B2(\RegFile/_3047_ ), .ZN(\RegFile/_0424_ ) );
AOI21_X1 \RegFile/_7459_ ( .A(\RegFile/_3793_ ), .B1(\RegFile/_3057_ ), .B2(\RegFile/_3058_ ), .ZN(\RegFile/_3061_ ) );
AOI21_X1 \RegFile/_7460_ ( .A(\RegFile/_3061_ ), .B1(\RegFile/_2299_ ), .B2(\RegFile/_3047_ ), .ZN(\RegFile/_0425_ ) );
NAND2_X1 \RegFile/_7461_ ( .A1(\RegFile/_3052_ ), .A2(\RegFile/_3763_ ), .ZN(\RegFile/_3062_ ) );
OAI21_X1 \RegFile/_7462_ ( .A(\RegFile/_3062_ ), .B1(\RegFile/_2317_ ), .B2(\RegFile/_3054_ ), .ZN(\RegFile/_0426_ ) );
AOI21_X1 \RegFile/_7463_ ( .A(\RegFile/_3764_ ), .B1(\RegFile/_3057_ ), .B2(\RegFile/_3058_ ), .ZN(\RegFile/_3063_ ) );
AOI21_X1 \RegFile/_7464_ ( .A(\RegFile/_3063_ ), .B1(\RegFile/_2336_ ), .B2(\RegFile/_3047_ ), .ZN(\RegFile/_0427_ ) );
AOI21_X1 \RegFile/_7465_ ( .A(\RegFile/_3765_ ), .B1(\RegFile/_3057_ ), .B2(\RegFile/_3058_ ), .ZN(\RegFile/_3064_ ) );
AOI21_X1 \RegFile/_7466_ ( .A(\RegFile/_3064_ ), .B1(\RegFile/_2356_ ), .B2(\RegFile/_3047_ ), .ZN(\RegFile/_0428_ ) );
AOI21_X1 \RegFile/_7467_ ( .A(\RegFile/_3766_ ), .B1(\RegFile/_3057_ ), .B2(\RegFile/_3058_ ), .ZN(\RegFile/_3065_ ) );
BUF_X4 \RegFile/_7468_ ( .A(\RegFile/_2014_ ), .Z(\RegFile/_3066_ ) );
AOI21_X1 \RegFile/_7469_ ( .A(\RegFile/_3065_ ), .B1(\RegFile/_2379_ ), .B2(\RegFile/_3066_ ), .ZN(\RegFile/_0429_ ) );
AOI21_X1 \RegFile/_7470_ ( .A(\RegFile/_3767_ ), .B1(\RegFile/_3057_ ), .B2(\RegFile/_3058_ ), .ZN(\RegFile/_3067_ ) );
AOI21_X1 \RegFile/_7471_ ( .A(\RegFile/_3067_ ), .B1(\RegFile/_2399_ ), .B2(\RegFile/_3066_ ), .ZN(\RegFile/_0430_ ) );
NAND2_X1 \RegFile/_7472_ ( .A1(\RegFile/_3052_ ), .A2(\RegFile/_3768_ ), .ZN(\RegFile/_3068_ ) );
OAI21_X1 \RegFile/_7473_ ( .A(\RegFile/_3068_ ), .B1(\RegFile/_2420_ ), .B2(\RegFile/_3054_ ), .ZN(\RegFile/_0431_ ) );
NAND2_X1 \RegFile/_7474_ ( .A1(\RegFile/_3052_ ), .A2(\RegFile/_3769_ ), .ZN(\RegFile/_3069_ ) );
OAI21_X1 \RegFile/_7475_ ( .A(\RegFile/_3069_ ), .B1(\RegFile/_2439_ ), .B2(\RegFile/_3054_ ), .ZN(\RegFile/_0432_ ) );
AOI21_X1 \RegFile/_7476_ ( .A(\RegFile/_3770_ ), .B1(\RegFile/_3057_ ), .B2(\RegFile/_3058_ ), .ZN(\RegFile/_3070_ ) );
AOI21_X1 \RegFile/_7477_ ( .A(\RegFile/_3070_ ), .B1(\RegFile/_2459_ ), .B2(\RegFile/_3066_ ), .ZN(\RegFile/_0433_ ) );
AOI21_X1 \RegFile/_7478_ ( .A(\RegFile/_3771_ ), .B1(\RegFile/_3057_ ), .B2(\RegFile/_3058_ ), .ZN(\RegFile/_3071_ ) );
AOI21_X1 \RegFile/_7479_ ( .A(\RegFile/_3071_ ), .B1(\RegFile/_2476_ ), .B2(\RegFile/_3066_ ), .ZN(\RegFile/_0434_ ) );
NAND2_X1 \RegFile/_7480_ ( .A1(\RegFile/_3052_ ), .A2(\RegFile/_3772_ ), .ZN(\RegFile/_3072_ ) );
OAI21_X1 \RegFile/_7481_ ( .A(\RegFile/_3072_ ), .B1(\RegFile/_2495_ ), .B2(\RegFile/_3054_ ), .ZN(\RegFile/_0435_ ) );
NAND2_X1 \RegFile/_7482_ ( .A1(\RegFile/_3052_ ), .A2(\RegFile/_3774_ ), .ZN(\RegFile/_3073_ ) );
OAI21_X1 \RegFile/_7483_ ( .A(\RegFile/_3073_ ), .B1(\RegFile/_2514_ ), .B2(\RegFile/_3054_ ), .ZN(\RegFile/_0436_ ) );
AOI21_X1 \RegFile/_7484_ ( .A(\RegFile/_3775_ ), .B1(\RegFile/_3057_ ), .B2(\RegFile/_3058_ ), .ZN(\RegFile/_3074_ ) );
AOI21_X1 \RegFile/_7485_ ( .A(\RegFile/_3074_ ), .B1(\RegFile/_2533_ ), .B2(\RegFile/_3066_ ), .ZN(\RegFile/_0437_ ) );
BUF_X4 \RegFile/_7486_ ( .A(\RegFile/_3006_ ), .Z(\RegFile/_3075_ ) );
AOI21_X1 \RegFile/_7487_ ( .A(\RegFile/_3776_ ), .B1(\RegFile/_3075_ ), .B2(\RegFile/_2725_ ), .ZN(\RegFile/_3076_ ) );
AOI21_X1 \RegFile/_7488_ ( .A(\RegFile/_3076_ ), .B1(\RegFile/_2552_ ), .B2(\RegFile/_3066_ ), .ZN(\RegFile/_0438_ ) );
AOI21_X1 \RegFile/_7489_ ( .A(\RegFile/_3777_ ), .B1(\RegFile/_3075_ ), .B2(\RegFile/_2725_ ), .ZN(\RegFile/_3077_ ) );
AOI21_X1 \RegFile/_7490_ ( .A(\RegFile/_3077_ ), .B1(\RegFile/_2571_ ), .B2(\RegFile/_3066_ ), .ZN(\RegFile/_0439_ ) );
AOI21_X1 \RegFile/_7491_ ( .A(\RegFile/_3778_ ), .B1(\RegFile/_3075_ ), .B2(\RegFile/_2725_ ), .ZN(\RegFile/_3078_ ) );
AOI21_X1 \RegFile/_7492_ ( .A(\RegFile/_3078_ ), .B1(\RegFile/_2592_ ), .B2(\RegFile/_3066_ ), .ZN(\RegFile/_0440_ ) );
AOI21_X1 \RegFile/_7493_ ( .A(\RegFile/_3779_ ), .B1(\RegFile/_3075_ ), .B2(\RegFile/_2725_ ), .ZN(\RegFile/_3079_ ) );
AOI21_X1 \RegFile/_7494_ ( .A(\RegFile/_3079_ ), .B1(\RegFile/_2608_ ), .B2(\RegFile/_3066_ ), .ZN(\RegFile/_0441_ ) );
NAND2_X1 \RegFile/_7495_ ( .A1(\RegFile/_3052_ ), .A2(\RegFile/_3780_ ), .ZN(\RegFile/_3080_ ) );
OAI21_X1 \RegFile/_7496_ ( .A(\RegFile/_3080_ ), .B1(\RegFile/_2627_ ), .B2(\RegFile/_3054_ ), .ZN(\RegFile/_0442_ ) );
AOI21_X1 \RegFile/_7497_ ( .A(\RegFile/_3781_ ), .B1(\RegFile/_3075_ ), .B2(\RegFile/_2725_ ), .ZN(\RegFile/_3081_ ) );
AOI21_X1 \RegFile/_7498_ ( .A(\RegFile/_3081_ ), .B1(\RegFile/_2646_ ), .B2(\RegFile/_3066_ ), .ZN(\RegFile/_0443_ ) );
NAND2_X1 \RegFile/_7499_ ( .A1(\RegFile/_3052_ ), .A2(\RegFile/_3782_ ), .ZN(\RegFile/_3082_ ) );
OAI21_X1 \RegFile/_7500_ ( .A(\RegFile/_3082_ ), .B1(\RegFile/_2664_ ), .B2(\RegFile/_3054_ ), .ZN(\RegFile/_0444_ ) );
NAND2_X1 \RegFile/_7501_ ( .A1(\RegFile/_3052_ ), .A2(\RegFile/_3783_ ), .ZN(\RegFile/_3083_ ) );
OAI21_X1 \RegFile/_7502_ ( .A(\RegFile/_3083_ ), .B1(\RegFile/_2684_ ), .B2(\RegFile/_3054_ ), .ZN(\RegFile/_0445_ ) );
AOI21_X1 \RegFile/_7503_ ( .A(\RegFile/_3785_ ), .B1(\RegFile/_3075_ ), .B2(\RegFile/_2725_ ), .ZN(\RegFile/_3084_ ) );
AOI21_X1 \RegFile/_7504_ ( .A(\RegFile/_3084_ ), .B1(\RegFile/_2705_ ), .B2(\RegFile/_2014_ ), .ZN(\RegFile/_0446_ ) );
AOI21_X1 \RegFile/_7505_ ( .A(\RegFile/_3786_ ), .B1(\RegFile/_3075_ ), .B2(\RegFile/_2725_ ), .ZN(\RegFile/_3085_ ) );
AOI21_X1 \RegFile/_7506_ ( .A(\RegFile/_3085_ ), .B1(\RegFile/_2724_ ), .B2(\RegFile/_2014_ ), .ZN(\RegFile/_0447_ ) );
INV_X1 \RegFile/_7507_ ( .A(\RegFile/_2206_ ), .ZN(\RegFile/_3086_ ) );
BUF_X4 \RegFile/_7508_ ( .A(\RegFile/_3086_ ), .Z(\RegFile/_3087_ ) );
NAND2_X1 \RegFile/_7509_ ( .A1(\RegFile/_3087_ ), .A2(\RegFile/_3314_ ), .ZN(\RegFile/_3088_ ) );
OAI21_X1 \RegFile/_7510_ ( .A(\RegFile/_3088_ ), .B1(\RegFile/_2071_ ), .B2(\RegFile/_3087_ ), .ZN(\RegFile/_0448_ ) );
NAND2_X1 \RegFile/_7511_ ( .A1(\RegFile/_3087_ ), .A2(\RegFile/_3325_ ), .ZN(\RegFile/_3089_ ) );
OAI21_X1 \RegFile/_7512_ ( .A(\RegFile/_3089_ ), .B1(\RegFile/_2113_ ), .B2(\RegFile/_3087_ ), .ZN(\RegFile/_0449_ ) );
AOI21_X1 \RegFile/_7513_ ( .A(\RegFile/_3336_ ), .B1(\RegFile/_3075_ ), .B2(\RegFile/_2802_ ), .ZN(\RegFile/_3090_ ) );
BUF_X4 \RegFile/_7514_ ( .A(\RegFile/_2206_ ), .Z(\RegFile/_3091_ ) );
AOI21_X1 \RegFile/_7515_ ( .A(\RegFile/_3090_ ), .B1(\RegFile/_2142_ ), .B2(\RegFile/_3091_ ), .ZN(\RegFile/_0450_ ) );
AOI21_X1 \RegFile/_7516_ ( .A(\RegFile/_3339_ ), .B1(\RegFile/_3075_ ), .B2(\RegFile/_2802_ ), .ZN(\RegFile/_3092_ ) );
AOI21_X1 \RegFile/_7517_ ( .A(\RegFile/_3092_ ), .B1(\RegFile/_2175_ ), .B2(\RegFile/_3091_ ), .ZN(\RegFile/_0451_ ) );
AOI21_X1 \RegFile/_7518_ ( .A(\RegFile/_3340_ ), .B1(\RegFile/_3075_ ), .B2(\RegFile/_2802_ ), .ZN(\RegFile/_3093_ ) );
AOI21_X1 \RegFile/_7519_ ( .A(\RegFile/_3093_ ), .B1(\RegFile/_2199_ ), .B2(\RegFile/_3091_ ), .ZN(\RegFile/_0452_ ) );
NAND2_X1 \RegFile/_7520_ ( .A1(\RegFile/_3087_ ), .A2(\RegFile/_3341_ ), .ZN(\RegFile/_3094_ ) );
OAI21_X1 \RegFile/_7521_ ( .A(\RegFile/_3094_ ), .B1(\RegFile/_2218_ ), .B2(\RegFile/_3087_ ), .ZN(\RegFile/_0453_ ) );
NAND2_X1 \RegFile/_7522_ ( .A1(\RegFile/_3086_ ), .A2(\RegFile/_3342_ ), .ZN(\RegFile/_3095_ ) );
OAI21_X1 \RegFile/_7523_ ( .A(\RegFile/_3095_ ), .B1(\RegFile/_2240_ ), .B2(\RegFile/_3087_ ), .ZN(\RegFile/_0454_ ) );
BUF_X4 \RegFile/_7524_ ( .A(\RegFile/_2160_ ), .Z(\RegFile/_3096_ ) );
AOI21_X1 \RegFile/_7525_ ( .A(\RegFile/_3343_ ), .B1(\RegFile/_3096_ ), .B2(\RegFile/_2802_ ), .ZN(\RegFile/_3097_ ) );
AOI21_X1 \RegFile/_7526_ ( .A(\RegFile/_3097_ ), .B1(\RegFile/_2261_ ), .B2(\RegFile/_3091_ ), .ZN(\RegFile/_0455_ ) );
AOI21_X1 \RegFile/_7527_ ( .A(\RegFile/_3344_ ), .B1(\RegFile/_3096_ ), .B2(\RegFile/_2802_ ), .ZN(\RegFile/_3098_ ) );
AOI21_X1 \RegFile/_7528_ ( .A(\RegFile/_3098_ ), .B1(\RegFile/_2782_ ), .B2(\RegFile/_3091_ ), .ZN(\RegFile/_0456_ ) );
AOI21_X1 \RegFile/_7529_ ( .A(\RegFile/_3345_ ), .B1(\RegFile/_3096_ ), .B2(\RegFile/_2802_ ), .ZN(\RegFile/_3099_ ) );
AOI21_X1 \RegFile/_7530_ ( .A(\RegFile/_3099_ ), .B1(\RegFile/_2299_ ), .B2(\RegFile/_3091_ ), .ZN(\RegFile/_0457_ ) );
AOI21_X1 \RegFile/_7531_ ( .A(\RegFile/_3315_ ), .B1(\RegFile/_3096_ ), .B2(\RegFile/_2802_ ), .ZN(\RegFile/_3100_ ) );
AOI21_X1 \RegFile/_7532_ ( .A(\RegFile/_3100_ ), .B1(\RegFile/_2318_ ), .B2(\RegFile/_3091_ ), .ZN(\RegFile/_0458_ ) );
BUF_X4 \RegFile/_7533_ ( .A(\RegFile/_2169_ ), .Z(\RegFile/_3101_ ) );
AOI21_X1 \RegFile/_7534_ ( .A(\RegFile/_3316_ ), .B1(\RegFile/_3096_ ), .B2(\RegFile/_3101_ ), .ZN(\RegFile/_3102_ ) );
AOI21_X1 \RegFile/_7535_ ( .A(\RegFile/_3102_ ), .B1(\RegFile/_2336_ ), .B2(\RegFile/_3091_ ), .ZN(\RegFile/_0459_ ) );
AOI21_X1 \RegFile/_7536_ ( .A(\RegFile/_3317_ ), .B1(\RegFile/_3096_ ), .B2(\RegFile/_3101_ ), .ZN(\RegFile/_3103_ ) );
AOI21_X1 \RegFile/_7537_ ( .A(\RegFile/_3103_ ), .B1(\RegFile/_2356_ ), .B2(\RegFile/_3091_ ), .ZN(\RegFile/_0460_ ) );
NAND2_X1 \RegFile/_7538_ ( .A1(\RegFile/_3086_ ), .A2(\RegFile/_3318_ ), .ZN(\RegFile/_3104_ ) );
OAI21_X1 \RegFile/_7539_ ( .A(\RegFile/_3104_ ), .B1(\RegFile/_2378_ ), .B2(\RegFile/_3087_ ), .ZN(\RegFile/_0461_ ) );
AOI21_X1 \RegFile/_7540_ ( .A(\RegFile/_3319_ ), .B1(\RegFile/_3096_ ), .B2(\RegFile/_3101_ ), .ZN(\RegFile/_3105_ ) );
AOI21_X1 \RegFile/_7541_ ( .A(\RegFile/_3105_ ), .B1(\RegFile/_2399_ ), .B2(\RegFile/_3091_ ), .ZN(\RegFile/_0462_ ) );
NAND2_X1 \RegFile/_7542_ ( .A1(\RegFile/_3086_ ), .A2(\RegFile/_3320_ ), .ZN(\RegFile/_3106_ ) );
OAI21_X1 \RegFile/_7543_ ( .A(\RegFile/_3106_ ), .B1(\RegFile/_2419_ ), .B2(\RegFile/_3087_ ), .ZN(\RegFile/_0463_ ) );
AOI21_X1 \RegFile/_7544_ ( .A(\RegFile/_3321_ ), .B1(\RegFile/_3096_ ), .B2(\RegFile/_3101_ ), .ZN(\RegFile/_3107_ ) );
BUF_X4 \RegFile/_7545_ ( .A(\RegFile/_2206_ ), .Z(\RegFile/_3108_ ) );
AOI21_X1 \RegFile/_7546_ ( .A(\RegFile/_3107_ ), .B1(\RegFile/_2440_ ), .B2(\RegFile/_3108_ ), .ZN(\RegFile/_0464_ ) );
AOI21_X1 \RegFile/_7547_ ( .A(\RegFile/_3322_ ), .B1(\RegFile/_3096_ ), .B2(\RegFile/_3101_ ), .ZN(\RegFile/_3109_ ) );
AOI21_X1 \RegFile/_7548_ ( .A(\RegFile/_3109_ ), .B1(\RegFile/_2459_ ), .B2(\RegFile/_3108_ ), .ZN(\RegFile/_0465_ ) );
AOI21_X1 \RegFile/_7549_ ( .A(\RegFile/_3323_ ), .B1(\RegFile/_3096_ ), .B2(\RegFile/_3101_ ), .ZN(\RegFile/_3110_ ) );
AOI21_X1 \RegFile/_7550_ ( .A(\RegFile/_3110_ ), .B1(\RegFile/_2476_ ), .B2(\RegFile/_3108_ ), .ZN(\RegFile/_0466_ ) );
BUF_X4 \RegFile/_7551_ ( .A(\RegFile/_2160_ ), .Z(\RegFile/_3111_ ) );
AOI21_X1 \RegFile/_7552_ ( .A(\RegFile/_3324_ ), .B1(\RegFile/_3111_ ), .B2(\RegFile/_3101_ ), .ZN(\RegFile/_3112_ ) );
AOI21_X1 \RegFile/_7553_ ( .A(\RegFile/_3112_ ), .B1(\RegFile/_2495_ ), .B2(\RegFile/_3108_ ), .ZN(\RegFile/_0467_ ) );
AOI21_X1 \RegFile/_7554_ ( .A(\RegFile/_3326_ ), .B1(\RegFile/_3111_ ), .B2(\RegFile/_3101_ ), .ZN(\RegFile/_3113_ ) );
AOI21_X1 \RegFile/_7555_ ( .A(\RegFile/_3113_ ), .B1(\RegFile/_2514_ ), .B2(\RegFile/_3108_ ), .ZN(\RegFile/_0468_ ) );
AOI21_X1 \RegFile/_7556_ ( .A(\RegFile/_3327_ ), .B1(\RegFile/_3111_ ), .B2(\RegFile/_3101_ ), .ZN(\RegFile/_3114_ ) );
AOI21_X1 \RegFile/_7557_ ( .A(\RegFile/_3114_ ), .B1(\RegFile/_2533_ ), .B2(\RegFile/_3108_ ), .ZN(\RegFile/_0469_ ) );
AOI21_X1 \RegFile/_7558_ ( .A(\RegFile/_3328_ ), .B1(\RegFile/_3111_ ), .B2(\RegFile/_3101_ ), .ZN(\RegFile/_3115_ ) );
AOI21_X1 \RegFile/_7559_ ( .A(\RegFile/_3115_ ), .B1(\RegFile/_2552_ ), .B2(\RegFile/_3108_ ), .ZN(\RegFile/_0470_ ) );
AOI21_X1 \RegFile/_7560_ ( .A(\RegFile/_3329_ ), .B1(\RegFile/_3111_ ), .B2(\RegFile/_2951_ ), .ZN(\RegFile/_3116_ ) );
AOI21_X1 \RegFile/_7561_ ( .A(\RegFile/_3116_ ), .B1(\RegFile/_2571_ ), .B2(\RegFile/_3108_ ), .ZN(\RegFile/_0471_ ) );
AOI21_X1 \RegFile/_7562_ ( .A(\RegFile/_3330_ ), .B1(\RegFile/_3111_ ), .B2(\RegFile/_2951_ ), .ZN(\RegFile/_3117_ ) );
AOI21_X1 \RegFile/_7563_ ( .A(\RegFile/_3117_ ), .B1(\RegFile/_2592_ ), .B2(\RegFile/_3108_ ), .ZN(\RegFile/_0472_ ) );
AOI21_X1 \RegFile/_7564_ ( .A(\RegFile/_3331_ ), .B1(\RegFile/_3111_ ), .B2(\RegFile/_2951_ ), .ZN(\RegFile/_3118_ ) );
AOI21_X1 \RegFile/_7565_ ( .A(\RegFile/_3118_ ), .B1(\RegFile/_2608_ ), .B2(\RegFile/_3108_ ), .ZN(\RegFile/_0473_ ) );
AOI21_X1 \RegFile/_7566_ ( .A(\RegFile/_3332_ ), .B1(\RegFile/_3111_ ), .B2(\RegFile/_2951_ ), .ZN(\RegFile/_3119_ ) );
AOI21_X1 \RegFile/_7567_ ( .A(\RegFile/_3119_ ), .B1(\RegFile/_2628_ ), .B2(\RegFile/_2206_ ), .ZN(\RegFile/_0474_ ) );
AOI21_X1 \RegFile/_7568_ ( .A(\RegFile/_3333_ ), .B1(\RegFile/_3111_ ), .B2(\RegFile/_2951_ ), .ZN(\RegFile/_3120_ ) );
AOI21_X1 \RegFile/_7569_ ( .A(\RegFile/_3120_ ), .B1(\RegFile/_2646_ ), .B2(\RegFile/_2206_ ), .ZN(\RegFile/_0475_ ) );
AOI21_X1 \RegFile/_7570_ ( .A(\RegFile/_3334_ ), .B1(\RegFile/_3111_ ), .B2(\RegFile/_2951_ ), .ZN(\RegFile/_3121_ ) );
AOI21_X1 \RegFile/_7571_ ( .A(\RegFile/_3121_ ), .B1(\RegFile/_2664_ ), .B2(\RegFile/_2206_ ), .ZN(\RegFile/_0476_ ) );
BUF_X4 \RegFile/_7572_ ( .A(\RegFile/_2160_ ), .Z(\RegFile/_3122_ ) );
AOI21_X1 \RegFile/_7573_ ( .A(\RegFile/_3335_ ), .B1(\RegFile/_3122_ ), .B2(\RegFile/_2951_ ), .ZN(\RegFile/_3123_ ) );
AOI21_X1 \RegFile/_7574_ ( .A(\RegFile/_3123_ ), .B1(\RegFile/_2685_ ), .B2(\RegFile/_2206_ ), .ZN(\RegFile/_0477_ ) );
NAND2_X1 \RegFile/_7575_ ( .A1(\RegFile/_3086_ ), .A2(\RegFile/_3337_ ), .ZN(\RegFile/_3124_ ) );
OAI21_X1 \RegFile/_7576_ ( .A(\RegFile/_3124_ ), .B1(\RegFile/_2704_ ), .B2(\RegFile/_3087_ ), .ZN(\RegFile/_0478_ ) );
AOI21_X1 \RegFile/_7577_ ( .A(\RegFile/_3338_ ), .B1(\RegFile/_3122_ ), .B2(\RegFile/_2951_ ), .ZN(\RegFile/_3125_ ) );
AOI21_X1 \RegFile/_7578_ ( .A(\RegFile/_3125_ ), .B1(\RegFile/_2724_ ), .B2(\RegFile/_2206_ ), .ZN(\RegFile/_0479_ ) );
AOI21_X1 \RegFile/_7579_ ( .A(\RegFile/_3346_ ), .B1(\RegFile/_3122_ ), .B2(\RegFile/_2839_ ), .ZN(\RegFile/_3126_ ) );
BUF_X4 \RegFile/_7580_ ( .A(\RegFile/_2021_ ), .Z(\RegFile/_3127_ ) );
AOI21_X1 \RegFile/_7581_ ( .A(\RegFile/_3126_ ), .B1(\RegFile/_2072_ ), .B2(\RegFile/_3127_ ), .ZN(\RegFile/_0480_ ) );
AOI21_X1 \RegFile/_7582_ ( .A(\RegFile/_3357_ ), .B1(\RegFile/_3122_ ), .B2(\RegFile/_2839_ ), .ZN(\RegFile/_3128_ ) );
AOI21_X1 \RegFile/_7583_ ( .A(\RegFile/_3128_ ), .B1(\RegFile/_2113_ ), .B2(\RegFile/_3127_ ), .ZN(\RegFile/_0481_ ) );
BUF_X4 \RegFile/_7584_ ( .A(\RegFile/_1990_ ), .Z(\RegFile/_3129_ ) );
AOI21_X1 \RegFile/_7585_ ( .A(\RegFile/_3368_ ), .B1(\RegFile/_3122_ ), .B2(\RegFile/_3129_ ), .ZN(\RegFile/_3130_ ) );
AOI21_X1 \RegFile/_7586_ ( .A(\RegFile/_3130_ ), .B1(\RegFile/_2142_ ), .B2(\RegFile/_3127_ ), .ZN(\RegFile/_0482_ ) );
AOI21_X1 \RegFile/_7587_ ( .A(\RegFile/_3371_ ), .B1(\RegFile/_3122_ ), .B2(\RegFile/_3129_ ), .ZN(\RegFile/_3131_ ) );
AOI21_X1 \RegFile/_7588_ ( .A(\RegFile/_3131_ ), .B1(\RegFile/_2175_ ), .B2(\RegFile/_3127_ ), .ZN(\RegFile/_0483_ ) );
AOI21_X1 \RegFile/_7589_ ( .A(\RegFile/_3372_ ), .B1(\RegFile/_3122_ ), .B2(\RegFile/_3129_ ), .ZN(\RegFile/_3132_ ) );
AOI21_X1 \RegFile/_7590_ ( .A(\RegFile/_3132_ ), .B1(\RegFile/_2199_ ), .B2(\RegFile/_3127_ ), .ZN(\RegFile/_0484_ ) );
INV_X2 \RegFile/_7591_ ( .A(\RegFile/_2021_ ), .ZN(\RegFile/_3133_ ) );
BUF_X4 \RegFile/_7592_ ( .A(\RegFile/_3133_ ), .Z(\RegFile/_3134_ ) );
NAND2_X1 \RegFile/_7593_ ( .A1(\RegFile/_3134_ ), .A2(\RegFile/_3373_ ), .ZN(\RegFile/_3135_ ) );
OAI21_X1 \RegFile/_7594_ ( .A(\RegFile/_3135_ ), .B1(\RegFile/_2218_ ), .B2(\RegFile/_3134_ ), .ZN(\RegFile/_0485_ ) );
AOI21_X1 \RegFile/_7595_ ( .A(\RegFile/_3374_ ), .B1(\RegFile/_3122_ ), .B2(\RegFile/_3129_ ), .ZN(\RegFile/_3136_ ) );
AOI21_X1 \RegFile/_7596_ ( .A(\RegFile/_3136_ ), .B1(\RegFile/_2240_ ), .B2(\RegFile/_3127_ ), .ZN(\RegFile/_0486_ ) );
AOI21_X1 \RegFile/_7597_ ( .A(\RegFile/_3375_ ), .B1(\RegFile/_3122_ ), .B2(\RegFile/_3129_ ), .ZN(\RegFile/_3137_ ) );
AOI21_X1 \RegFile/_7598_ ( .A(\RegFile/_3137_ ), .B1(\RegFile/_2261_ ), .B2(\RegFile/_3127_ ), .ZN(\RegFile/_0487_ ) );
AOI21_X1 \RegFile/_7599_ ( .A(\RegFile/_3376_ ), .B1(\RegFile/_3122_ ), .B2(\RegFile/_3129_ ), .ZN(\RegFile/_3138_ ) );
AOI21_X1 \RegFile/_7600_ ( .A(\RegFile/_3138_ ), .B1(\RegFile/_2782_ ), .B2(\RegFile/_3127_ ), .ZN(\RegFile/_0488_ ) );
BUF_X4 \RegFile/_7601_ ( .A(\RegFile/_2160_ ), .Z(\RegFile/_3139_ ) );
AOI21_X1 \RegFile/_7602_ ( .A(\RegFile/_3377_ ), .B1(\RegFile/_3139_ ), .B2(\RegFile/_3129_ ), .ZN(\RegFile/_3140_ ) );
AOI21_X1 \RegFile/_7603_ ( .A(\RegFile/_3140_ ), .B1(\RegFile/_2299_ ), .B2(\RegFile/_3127_ ), .ZN(\RegFile/_0489_ ) );
AOI21_X1 \RegFile/_7604_ ( .A(\RegFile/_3347_ ), .B1(\RegFile/_3139_ ), .B2(\RegFile/_3129_ ), .ZN(\RegFile/_3141_ ) );
AOI21_X1 \RegFile/_7605_ ( .A(\RegFile/_3141_ ), .B1(\RegFile/_2318_ ), .B2(\RegFile/_3127_ ), .ZN(\RegFile/_0490_ ) );
AOI21_X1 \RegFile/_7606_ ( .A(\RegFile/_3348_ ), .B1(\RegFile/_3139_ ), .B2(\RegFile/_3129_ ), .ZN(\RegFile/_3142_ ) );
BUF_X4 \RegFile/_7607_ ( .A(\RegFile/_2021_ ), .Z(\RegFile/_3143_ ) );
AOI21_X1 \RegFile/_7608_ ( .A(\RegFile/_3142_ ), .B1(\RegFile/_2336_ ), .B2(\RegFile/_3143_ ), .ZN(\RegFile/_0491_ ) );
AOI21_X1 \RegFile/_7609_ ( .A(\RegFile/_3349_ ), .B1(\RegFile/_3139_ ), .B2(\RegFile/_3129_ ), .ZN(\RegFile/_3144_ ) );
AOI21_X1 \RegFile/_7610_ ( .A(\RegFile/_3144_ ), .B1(\RegFile/_2356_ ), .B2(\RegFile/_3143_ ), .ZN(\RegFile/_0492_ ) );
BUF_X4 \RegFile/_7611_ ( .A(\RegFile/_1990_ ), .Z(\RegFile/_3145_ ) );
AOI21_X1 \RegFile/_7612_ ( .A(\RegFile/_3350_ ), .B1(\RegFile/_3139_ ), .B2(\RegFile/_3145_ ), .ZN(\RegFile/_3146_ ) );
AOI21_X1 \RegFile/_7613_ ( .A(\RegFile/_3146_ ), .B1(\RegFile/_2379_ ), .B2(\RegFile/_3143_ ), .ZN(\RegFile/_0493_ ) );
NAND2_X1 \RegFile/_7614_ ( .A1(\RegFile/_3133_ ), .A2(\RegFile/_3351_ ), .ZN(\RegFile/_3147_ ) );
OAI21_X1 \RegFile/_7615_ ( .A(\RegFile/_3147_ ), .B1(\RegFile/_2399_ ), .B2(\RegFile/_3134_ ), .ZN(\RegFile/_0494_ ) );
NAND2_X1 \RegFile/_7616_ ( .A1(\RegFile/_3133_ ), .A2(\RegFile/_3352_ ), .ZN(\RegFile/_3148_ ) );
OAI21_X1 \RegFile/_7617_ ( .A(\RegFile/_3148_ ), .B1(\RegFile/_2419_ ), .B2(\RegFile/_3134_ ), .ZN(\RegFile/_0495_ ) );
NAND2_X1 \RegFile/_7618_ ( .A1(\RegFile/_3133_ ), .A2(\RegFile/_3353_ ), .ZN(\RegFile/_3149_ ) );
OAI21_X1 \RegFile/_7619_ ( .A(\RegFile/_3149_ ), .B1(\RegFile/_2439_ ), .B2(\RegFile/_3134_ ), .ZN(\RegFile/_0496_ ) );
AOI21_X1 \RegFile/_7620_ ( .A(\RegFile/_3354_ ), .B1(\RegFile/_3139_ ), .B2(\RegFile/_3145_ ), .ZN(\RegFile/_3150_ ) );
AOI21_X1 \RegFile/_7621_ ( .A(\RegFile/_3150_ ), .B1(\RegFile/_2459_ ), .B2(\RegFile/_3143_ ), .ZN(\RegFile/_0497_ ) );
NAND2_X1 \RegFile/_7622_ ( .A1(\RegFile/_3133_ ), .A2(\RegFile/_3355_ ), .ZN(\RegFile/_3151_ ) );
OAI21_X1 \RegFile/_7623_ ( .A(\RegFile/_3151_ ), .B1(\RegFile/_2476_ ), .B2(\RegFile/_3134_ ), .ZN(\RegFile/_0498_ ) );
AOI21_X1 \RegFile/_7624_ ( .A(\RegFile/_3356_ ), .B1(\RegFile/_3139_ ), .B2(\RegFile/_3145_ ), .ZN(\RegFile/_3152_ ) );
AOI21_X1 \RegFile/_7625_ ( .A(\RegFile/_3152_ ), .B1(\RegFile/_2495_ ), .B2(\RegFile/_3143_ ), .ZN(\RegFile/_0499_ ) );
AOI21_X1 \RegFile/_7626_ ( .A(\RegFile/_3358_ ), .B1(\RegFile/_3139_ ), .B2(\RegFile/_3145_ ), .ZN(\RegFile/_3153_ ) );
AOI21_X1 \RegFile/_7627_ ( .A(\RegFile/_3153_ ), .B1(\RegFile/_2514_ ), .B2(\RegFile/_3143_ ), .ZN(\RegFile/_0500_ ) );
NAND2_X1 \RegFile/_7628_ ( .A1(\RegFile/_3133_ ), .A2(\RegFile/_3359_ ), .ZN(\RegFile/_3154_ ) );
OAI21_X1 \RegFile/_7629_ ( .A(\RegFile/_3154_ ), .B1(\RegFile/_2533_ ), .B2(\RegFile/_3134_ ), .ZN(\RegFile/_0501_ ) );
AOI21_X1 \RegFile/_7630_ ( .A(\RegFile/_3360_ ), .B1(\RegFile/_3139_ ), .B2(\RegFile/_3145_ ), .ZN(\RegFile/_3155_ ) );
AOI21_X1 \RegFile/_7631_ ( .A(\RegFile/_3155_ ), .B1(\RegFile/_2552_ ), .B2(\RegFile/_3143_ ), .ZN(\RegFile/_0502_ ) );
NAND2_X1 \RegFile/_7632_ ( .A1(\RegFile/_3133_ ), .A2(\RegFile/_3361_ ), .ZN(\RegFile/_3156_ ) );
OAI21_X1 \RegFile/_7633_ ( .A(\RegFile/_3156_ ), .B1(\RegFile/_2571_ ), .B2(\RegFile/_3134_ ), .ZN(\RegFile/_0503_ ) );
NAND2_X1 \RegFile/_7634_ ( .A1(\RegFile/_3133_ ), .A2(\RegFile/_3362_ ), .ZN(\RegFile/_3157_ ) );
OAI21_X1 \RegFile/_7635_ ( .A(\RegFile/_3157_ ), .B1(\RegFile/_2591_ ), .B2(\RegFile/_3134_ ), .ZN(\RegFile/_0504_ ) );
AOI21_X1 \RegFile/_7636_ ( .A(\RegFile/_3363_ ), .B1(\RegFile/_3139_ ), .B2(\RegFile/_3145_ ), .ZN(\RegFile/_3158_ ) );
AOI21_X1 \RegFile/_7637_ ( .A(\RegFile/_3158_ ), .B1(\RegFile/_2608_ ), .B2(\RegFile/_3143_ ), .ZN(\RegFile/_0505_ ) );
AOI21_X1 \RegFile/_7638_ ( .A(\RegFile/_3364_ ), .B1(\RegFile/_3006_ ), .B2(\RegFile/_3145_ ), .ZN(\RegFile/_3159_ ) );
AOI21_X1 \RegFile/_7639_ ( .A(\RegFile/_3159_ ), .B1(\RegFile/_2628_ ), .B2(\RegFile/_3143_ ), .ZN(\RegFile/_0506_ ) );
AOI21_X1 \RegFile/_7640_ ( .A(\RegFile/_3365_ ), .B1(\RegFile/_3006_ ), .B2(\RegFile/_3145_ ), .ZN(\RegFile/_3160_ ) );
AOI21_X1 \RegFile/_7641_ ( .A(\RegFile/_3160_ ), .B1(\RegFile/_2646_ ), .B2(\RegFile/_3143_ ), .ZN(\RegFile/_0507_ ) );
NAND2_X1 \RegFile/_7642_ ( .A1(\RegFile/_3133_ ), .A2(\RegFile/_3366_ ), .ZN(\RegFile/_3161_ ) );
OAI21_X1 \RegFile/_7643_ ( .A(\RegFile/_3161_ ), .B1(\RegFile/_2663_ ), .B2(\RegFile/_3134_ ), .ZN(\RegFile/_0508_ ) );
AOI21_X1 \RegFile/_7644_ ( .A(\RegFile/_3367_ ), .B1(\RegFile/_3006_ ), .B2(\RegFile/_3145_ ), .ZN(\RegFile/_3162_ ) );
AOI21_X1 \RegFile/_7645_ ( .A(\RegFile/_3162_ ), .B1(\RegFile/_2685_ ), .B2(\RegFile/_2021_ ), .ZN(\RegFile/_0509_ ) );
AOI21_X1 \RegFile/_7646_ ( .A(\RegFile/_3369_ ), .B1(\RegFile/_3006_ ), .B2(\RegFile/_3145_ ), .ZN(\RegFile/_3163_ ) );
AOI21_X1 \RegFile/_7647_ ( .A(\RegFile/_3163_ ), .B1(\RegFile/_2705_ ), .B2(\RegFile/_2021_ ), .ZN(\RegFile/_0510_ ) );
AOI21_X1 \RegFile/_7648_ ( .A(\RegFile/_3370_ ), .B1(\RegFile/_3006_ ), .B2(\RegFile/_1990_ ), .ZN(\RegFile/_3164_ ) );
AOI21_X1 \RegFile/_7649_ ( .A(\RegFile/_3164_ ), .B1(\RegFile/_2724_ ), .B2(\RegFile/_2021_ ), .ZN(\RegFile/_0511_ ) );
BUF_X4 \RegFile/_7650_ ( .A(\RegFile/_1996_ ), .Z(\RegFile/_3165_ ) );
BUF_X4 \RegFile/_7651_ ( .A(\RegFile/_3165_ ), .Z(\RegFile/_3166_ ) );
AOI21_X1 \RegFile/_7652_ ( .A(\RegFile/_3378_ ), .B1(\RegFile/_3166_ ), .B2(\RegFile/_3035_ ), .ZN(\RegFile/_3167_ ) );
BUF_X4 \RegFile/_7653_ ( .A(\RegFile/_2024_ ), .Z(\RegFile/_3168_ ) );
AOI21_X1 \RegFile/_7654_ ( .A(\RegFile/_3167_ ), .B1(\RegFile/_2072_ ), .B2(\RegFile/_3168_ ), .ZN(\RegFile/_0512_ ) );
INV_X1 \RegFile/_7655_ ( .A(\RegFile/_2024_ ), .ZN(\RegFile/_3169_ ) );
BUF_X4 \RegFile/_7656_ ( .A(\RegFile/_3169_ ), .Z(\RegFile/_3170_ ) );
NAND2_X1 \RegFile/_7657_ ( .A1(\RegFile/_3170_ ), .A2(\RegFile/_3389_ ), .ZN(\RegFile/_3171_ ) );
BUF_X4 \RegFile/_7658_ ( .A(\RegFile/_3169_ ), .Z(\RegFile/_3172_ ) );
OAI21_X1 \RegFile/_7659_ ( .A(\RegFile/_3171_ ), .B1(\RegFile/_2113_ ), .B2(\RegFile/_3172_ ), .ZN(\RegFile/_0513_ ) );
AOI21_X1 \RegFile/_7660_ ( .A(\RegFile/_3400_ ), .B1(\RegFile/_3166_ ), .B2(\RegFile/_3035_ ), .ZN(\RegFile/_3173_ ) );
AOI21_X1 \RegFile/_7661_ ( .A(\RegFile/_3173_ ), .B1(\RegFile/_2142_ ), .B2(\RegFile/_3168_ ), .ZN(\RegFile/_0514_ ) );
AOI21_X1 \RegFile/_7662_ ( .A(\RegFile/_3403_ ), .B1(\RegFile/_3166_ ), .B2(\RegFile/_3035_ ), .ZN(\RegFile/_3174_ ) );
AOI21_X1 \RegFile/_7663_ ( .A(\RegFile/_3174_ ), .B1(\RegFile/_2175_ ), .B2(\RegFile/_3168_ ), .ZN(\RegFile/_0515_ ) );
BUF_X4 \RegFile/_7664_ ( .A(\RegFile/_2035_ ), .Z(\RegFile/_3175_ ) );
AOI21_X1 \RegFile/_7665_ ( .A(\RegFile/_3404_ ), .B1(\RegFile/_3166_ ), .B2(\RegFile/_3175_ ), .ZN(\RegFile/_3176_ ) );
AOI21_X1 \RegFile/_7666_ ( .A(\RegFile/_3176_ ), .B1(\RegFile/_2199_ ), .B2(\RegFile/_3168_ ), .ZN(\RegFile/_0516_ ) );
NAND2_X1 \RegFile/_7667_ ( .A1(\RegFile/_3170_ ), .A2(\RegFile/_3405_ ), .ZN(\RegFile/_3177_ ) );
OAI21_X1 \RegFile/_7668_ ( .A(\RegFile/_3177_ ), .B1(\RegFile/_2218_ ), .B2(\RegFile/_3172_ ), .ZN(\RegFile/_0517_ ) );
NAND2_X1 \RegFile/_7669_ ( .A1(\RegFile/_3170_ ), .A2(\RegFile/_3406_ ), .ZN(\RegFile/_3178_ ) );
OAI21_X1 \RegFile/_7670_ ( .A(\RegFile/_3178_ ), .B1(\RegFile/_2239_ ), .B2(\RegFile/_3172_ ), .ZN(\RegFile/_0518_ ) );
AOI21_X1 \RegFile/_7671_ ( .A(\RegFile/_3407_ ), .B1(\RegFile/_3166_ ), .B2(\RegFile/_3175_ ), .ZN(\RegFile/_3179_ ) );
AOI21_X1 \RegFile/_7672_ ( .A(\RegFile/_3179_ ), .B1(\RegFile/_2261_ ), .B2(\RegFile/_3168_ ), .ZN(\RegFile/_0519_ ) );
AOI21_X1 \RegFile/_7673_ ( .A(\RegFile/_3408_ ), .B1(\RegFile/_3166_ ), .B2(\RegFile/_3175_ ), .ZN(\RegFile/_3180_ ) );
AOI21_X1 \RegFile/_7674_ ( .A(\RegFile/_3180_ ), .B1(\RegFile/_2782_ ), .B2(\RegFile/_3168_ ), .ZN(\RegFile/_0520_ ) );
NAND2_X1 \RegFile/_7675_ ( .A1(\RegFile/_3170_ ), .A2(\RegFile/_3409_ ), .ZN(\RegFile/_3181_ ) );
OAI21_X1 \RegFile/_7676_ ( .A(\RegFile/_3181_ ), .B1(\RegFile/_2299_ ), .B2(\RegFile/_3172_ ), .ZN(\RegFile/_0521_ ) );
AOI21_X1 \RegFile/_7677_ ( .A(\RegFile/_3379_ ), .B1(\RegFile/_3166_ ), .B2(\RegFile/_3175_ ), .ZN(\RegFile/_3182_ ) );
AOI21_X1 \RegFile/_7678_ ( .A(\RegFile/_3182_ ), .B1(\RegFile/_2318_ ), .B2(\RegFile/_3168_ ), .ZN(\RegFile/_0522_ ) );
NAND2_X1 \RegFile/_7679_ ( .A1(\RegFile/_3170_ ), .A2(\RegFile/_3380_ ), .ZN(\RegFile/_3183_ ) );
OAI21_X1 \RegFile/_7680_ ( .A(\RegFile/_3183_ ), .B1(\RegFile/_2336_ ), .B2(\RegFile/_3172_ ), .ZN(\RegFile/_0523_ ) );
AOI21_X1 \RegFile/_7681_ ( .A(\RegFile/_3381_ ), .B1(\RegFile/_3166_ ), .B2(\RegFile/_3175_ ), .ZN(\RegFile/_3184_ ) );
AOI21_X1 \RegFile/_7682_ ( .A(\RegFile/_3184_ ), .B1(\RegFile/_2356_ ), .B2(\RegFile/_3168_ ), .ZN(\RegFile/_0524_ ) );
AOI21_X1 \RegFile/_7683_ ( .A(\RegFile/_3382_ ), .B1(\RegFile/_3166_ ), .B2(\RegFile/_3175_ ), .ZN(\RegFile/_3185_ ) );
AOI21_X1 \RegFile/_7684_ ( .A(\RegFile/_3185_ ), .B1(\RegFile/_2379_ ), .B2(\RegFile/_3168_ ), .ZN(\RegFile/_0525_ ) );
AOI21_X1 \RegFile/_7685_ ( .A(\RegFile/_3383_ ), .B1(\RegFile/_3166_ ), .B2(\RegFile/_3175_ ), .ZN(\RegFile/_3186_ ) );
AOI21_X1 \RegFile/_7686_ ( .A(\RegFile/_3186_ ), .B1(\RegFile/_2399_ ), .B2(\RegFile/_3168_ ), .ZN(\RegFile/_0526_ ) );
BUF_X4 \RegFile/_7687_ ( .A(\RegFile/_3165_ ), .Z(\RegFile/_3187_ ) );
AOI21_X1 \RegFile/_7688_ ( .A(\RegFile/_3384_ ), .B1(\RegFile/_3187_ ), .B2(\RegFile/_3175_ ), .ZN(\RegFile/_3188_ ) );
BUF_X4 \RegFile/_7689_ ( .A(\RegFile/_2024_ ), .Z(\RegFile/_3189_ ) );
AOI21_X1 \RegFile/_7690_ ( .A(\RegFile/_3188_ ), .B1(\RegFile/_2420_ ), .B2(\RegFile/_3189_ ), .ZN(\RegFile/_0527_ ) );
AOI21_X1 \RegFile/_7691_ ( .A(\RegFile/_3385_ ), .B1(\RegFile/_3187_ ), .B2(\RegFile/_3175_ ), .ZN(\RegFile/_3190_ ) );
AOI21_X1 \RegFile/_7692_ ( .A(\RegFile/_3190_ ), .B1(\RegFile/_2440_ ), .B2(\RegFile/_3189_ ), .ZN(\RegFile/_0528_ ) );
AOI21_X1 \RegFile/_7693_ ( .A(\RegFile/_3386_ ), .B1(\RegFile/_3187_ ), .B2(\RegFile/_3175_ ), .ZN(\RegFile/_3191_ ) );
AOI21_X1 \RegFile/_7694_ ( .A(\RegFile/_3191_ ), .B1(\RegFile/_2459_ ), .B2(\RegFile/_3189_ ), .ZN(\RegFile/_0529_ ) );
AOI21_X1 \RegFile/_7695_ ( .A(\RegFile/_3387_ ), .B1(\RegFile/_3187_ ), .B2(\RegFile/_2847_ ), .ZN(\RegFile/_3192_ ) );
AOI21_X1 \RegFile/_7696_ ( .A(\RegFile/_3192_ ), .B1(\RegFile/_2476_ ), .B2(\RegFile/_3189_ ), .ZN(\RegFile/_0530_ ) );
NAND2_X1 \RegFile/_7697_ ( .A1(\RegFile/_3170_ ), .A2(\RegFile/_3388_ ), .ZN(\RegFile/_3193_ ) );
OAI21_X1 \RegFile/_7698_ ( .A(\RegFile/_3193_ ), .B1(\RegFile/_2495_ ), .B2(\RegFile/_3172_ ), .ZN(\RegFile/_0531_ ) );
AOI21_X1 \RegFile/_7699_ ( .A(\RegFile/_3390_ ), .B1(\RegFile/_3187_ ), .B2(\RegFile/_2847_ ), .ZN(\RegFile/_3194_ ) );
AOI21_X1 \RegFile/_7700_ ( .A(\RegFile/_3194_ ), .B1(\RegFile/_2514_ ), .B2(\RegFile/_3189_ ), .ZN(\RegFile/_0532_ ) );
NAND2_X1 \RegFile/_7701_ ( .A1(\RegFile/_3170_ ), .A2(\RegFile/_3391_ ), .ZN(\RegFile/_3195_ ) );
OAI21_X1 \RegFile/_7702_ ( .A(\RegFile/_3195_ ), .B1(\RegFile/_2533_ ), .B2(\RegFile/_3172_ ), .ZN(\RegFile/_0533_ ) );
NAND2_X1 \RegFile/_7703_ ( .A1(\RegFile/_3170_ ), .A2(\RegFile/_3392_ ), .ZN(\RegFile/_3196_ ) );
OAI21_X1 \RegFile/_7704_ ( .A(\RegFile/_3196_ ), .B1(\RegFile/_2552_ ), .B2(\RegFile/_3172_ ), .ZN(\RegFile/_0534_ ) );
NAND2_X1 \RegFile/_7705_ ( .A1(\RegFile/_3170_ ), .A2(\RegFile/_3393_ ), .ZN(\RegFile/_3197_ ) );
OAI21_X1 \RegFile/_7706_ ( .A(\RegFile/_3197_ ), .B1(\RegFile/_2571_ ), .B2(\RegFile/_3172_ ), .ZN(\RegFile/_0535_ ) );
NAND2_X1 \RegFile/_7707_ ( .A1(\RegFile/_3169_ ), .A2(\RegFile/_3394_ ), .ZN(\RegFile/_3198_ ) );
OAI21_X1 \RegFile/_7708_ ( .A(\RegFile/_3198_ ), .B1(\RegFile/_2591_ ), .B2(\RegFile/_3172_ ), .ZN(\RegFile/_0536_ ) );
NAND2_X1 \RegFile/_7709_ ( .A1(\RegFile/_3169_ ), .A2(\RegFile/_3395_ ), .ZN(\RegFile/_3199_ ) );
OAI21_X1 \RegFile/_7710_ ( .A(\RegFile/_3199_ ), .B1(\RegFile/_2608_ ), .B2(\RegFile/_3170_ ), .ZN(\RegFile/_0537_ ) );
AOI21_X1 \RegFile/_7711_ ( .A(\RegFile/_3396_ ), .B1(\RegFile/_3187_ ), .B2(\RegFile/_2847_ ), .ZN(\RegFile/_3200_ ) );
AOI21_X1 \RegFile/_7712_ ( .A(\RegFile/_3200_ ), .B1(\RegFile/_2628_ ), .B2(\RegFile/_3189_ ), .ZN(\RegFile/_0538_ ) );
AOI21_X1 \RegFile/_7713_ ( .A(\RegFile/_3397_ ), .B1(\RegFile/_3187_ ), .B2(\RegFile/_2847_ ), .ZN(\RegFile/_3201_ ) );
AOI21_X1 \RegFile/_7714_ ( .A(\RegFile/_3201_ ), .B1(\RegFile/_2646_ ), .B2(\RegFile/_3189_ ), .ZN(\RegFile/_0539_ ) );
AOI21_X1 \RegFile/_7715_ ( .A(\RegFile/_3398_ ), .B1(\RegFile/_3187_ ), .B2(\RegFile/_2847_ ), .ZN(\RegFile/_3202_ ) );
AOI21_X1 \RegFile/_7716_ ( .A(\RegFile/_3202_ ), .B1(\RegFile/_2664_ ), .B2(\RegFile/_3189_ ), .ZN(\RegFile/_0540_ ) );
AOI21_X1 \RegFile/_7717_ ( .A(\RegFile/_3399_ ), .B1(\RegFile/_3187_ ), .B2(\RegFile/_2847_ ), .ZN(\RegFile/_3203_ ) );
AOI21_X1 \RegFile/_7718_ ( .A(\RegFile/_3203_ ), .B1(\RegFile/_2685_ ), .B2(\RegFile/_3189_ ), .ZN(\RegFile/_0541_ ) );
AOI21_X1 \RegFile/_7719_ ( .A(\RegFile/_3401_ ), .B1(\RegFile/_3187_ ), .B2(\RegFile/_2847_ ), .ZN(\RegFile/_3204_ ) );
AOI21_X1 \RegFile/_7720_ ( .A(\RegFile/_3204_ ), .B1(\RegFile/_2705_ ), .B2(\RegFile/_3189_ ), .ZN(\RegFile/_0542_ ) );
AOI21_X1 \RegFile/_7721_ ( .A(\RegFile/_3402_ ), .B1(\RegFile/_1997_ ), .B2(\RegFile/_2847_ ), .ZN(\RegFile/_3205_ ) );
AOI21_X1 \RegFile/_7722_ ( .A(\RegFile/_3205_ ), .B1(\RegFile/_2724_ ), .B2(\RegFile/_2024_ ), .ZN(\RegFile/_0543_ ) );
AOI21_X1 \RegFile/_7723_ ( .A(\RegFile/_3410_ ), .B1(\RegFile/_2898_ ), .B2(\RegFile/_2665_ ), .ZN(\RegFile/_3206_ ) );
BUF_X4 \RegFile/_7724_ ( .A(\RegFile/_2031_ ), .Z(\RegFile/_3207_ ) );
AOI21_X1 \RegFile/_7725_ ( .A(\RegFile/_3206_ ), .B1(\RegFile/_2072_ ), .B2(\RegFile/_3207_ ), .ZN(\RegFile/_0544_ ) );
AOI21_X1 \RegFile/_7726_ ( .A(\RegFile/_2404_ ), .B1(\RegFile/_2110_ ), .B2(\RegFile/_2111_ ), .ZN(\RegFile/_3208_ ) );
BUF_X4 \RegFile/_7727_ ( .A(\RegFile/_2404_ ), .Z(\RegFile/_3209_ ) );
AOI21_X1 \RegFile/_7728_ ( .A(\RegFile/_3208_ ), .B1(\RegFile/_1459_ ), .B2(\RegFile/_3209_ ), .ZN(\RegFile/_0545_ ) );
BUF_X4 \RegFile/_7729_ ( .A(\RegFile/_2161_ ), .Z(\RegFile/_3210_ ) );
AOI21_X1 \RegFile/_7730_ ( .A(\RegFile/_3432_ ), .B1(\RegFile/_3210_ ), .B2(\RegFile/_2665_ ), .ZN(\RegFile/_3211_ ) );
AOI21_X1 \RegFile/_7731_ ( .A(\RegFile/_3211_ ), .B1(\RegFile/_2142_ ), .B2(\RegFile/_3207_ ), .ZN(\RegFile/_0546_ ) );
BUF_X4 \RegFile/_7732_ ( .A(\RegFile/_2404_ ), .Z(\RegFile/_3212_ ) );
NAND2_X1 \RegFile/_7733_ ( .A1(\RegFile/_3212_ ), .A2(\RegFile/_3435_ ), .ZN(\RegFile/_3213_ ) );
OAI21_X1 \RegFile/_7734_ ( .A(\RegFile/_3213_ ), .B1(\RegFile/_2175_ ), .B2(\RegFile/_3209_ ), .ZN(\RegFile/_0547_ ) );
NAND2_X1 \RegFile/_7735_ ( .A1(\RegFile/_3212_ ), .A2(\RegFile/_3436_ ), .ZN(\RegFile/_3214_ ) );
OAI21_X1 \RegFile/_7736_ ( .A(\RegFile/_3214_ ), .B1(\RegFile/_2199_ ), .B2(\RegFile/_3209_ ), .ZN(\RegFile/_0548_ ) );
AOI21_X1 \RegFile/_7737_ ( .A(\RegFile/_3437_ ), .B1(\RegFile/_3210_ ), .B2(\RegFile/_2665_ ), .ZN(\RegFile/_3215_ ) );
AOI21_X1 \RegFile/_7738_ ( .A(\RegFile/_3215_ ), .B1(\RegFile/_2218_ ), .B2(\RegFile/_3207_ ), .ZN(\RegFile/_0549_ ) );
AOI21_X1 \RegFile/_7739_ ( .A(\RegFile/_3438_ ), .B1(\RegFile/_3210_ ), .B2(\RegFile/_2665_ ), .ZN(\RegFile/_3216_ ) );
AOI21_X1 \RegFile/_7740_ ( .A(\RegFile/_3216_ ), .B1(\RegFile/_2240_ ), .B2(\RegFile/_3207_ ), .ZN(\RegFile/_0550_ ) );
AOI21_X1 \RegFile/_7741_ ( .A(\RegFile/_3439_ ), .B1(\RegFile/_3210_ ), .B2(\RegFile/_2665_ ), .ZN(\RegFile/_3217_ ) );
AOI21_X1 \RegFile/_7742_ ( .A(\RegFile/_3217_ ), .B1(\RegFile/_2261_ ), .B2(\RegFile/_3207_ ), .ZN(\RegFile/_0551_ ) );
AOI21_X1 \RegFile/_7743_ ( .A(\RegFile/_3440_ ), .B1(\RegFile/_3210_ ), .B2(\RegFile/_2665_ ), .ZN(\RegFile/_3218_ ) );
AOI21_X1 \RegFile/_7744_ ( .A(\RegFile/_3218_ ), .B1(\RegFile/_2782_ ), .B2(\RegFile/_3207_ ), .ZN(\RegFile/_0552_ ) );
NAND2_X1 \RegFile/_7745_ ( .A1(\RegFile/_3212_ ), .A2(\RegFile/_3441_ ), .ZN(\RegFile/_3219_ ) );
OAI21_X1 \RegFile/_7746_ ( .A(\RegFile/_3219_ ), .B1(\RegFile/_2299_ ), .B2(\RegFile/_3209_ ), .ZN(\RegFile/_0553_ ) );
AOI21_X1 \RegFile/_7747_ ( .A(\RegFile/_3411_ ), .B1(\RegFile/_3210_ ), .B2(\RegFile/_2665_ ), .ZN(\RegFile/_3220_ ) );
AOI21_X1 \RegFile/_7748_ ( .A(\RegFile/_3220_ ), .B1(\RegFile/_2318_ ), .B2(\RegFile/_3207_ ), .ZN(\RegFile/_0554_ ) );
AOI21_X1 \RegFile/_7749_ ( .A(\RegFile/_3412_ ), .B1(\RegFile/_3210_ ), .B2(\RegFile/_2665_ ), .ZN(\RegFile/_3221_ ) );
AOI21_X1 \RegFile/_7750_ ( .A(\RegFile/_3221_ ), .B1(\RegFile/_2336_ ), .B2(\RegFile/_3207_ ), .ZN(\RegFile/_0555_ ) );
AOI21_X1 \RegFile/_7751_ ( .A(\RegFile/_3413_ ), .B1(\RegFile/_3210_ ), .B2(\RegFile/_3165_ ), .ZN(\RegFile/_3222_ ) );
AOI21_X1 \RegFile/_7752_ ( .A(\RegFile/_3222_ ), .B1(\RegFile/_2356_ ), .B2(\RegFile/_3207_ ), .ZN(\RegFile/_0556_ ) );
NAND2_X1 \RegFile/_7753_ ( .A1(\RegFile/_3212_ ), .A2(\RegFile/_3414_ ), .ZN(\RegFile/_3223_ ) );
OAI21_X1 \RegFile/_7754_ ( .A(\RegFile/_3223_ ), .B1(\RegFile/_2378_ ), .B2(\RegFile/_3209_ ), .ZN(\RegFile/_0557_ ) );
NAND2_X1 \RegFile/_7755_ ( .A1(\RegFile/_3212_ ), .A2(\RegFile/_3415_ ), .ZN(\RegFile/_3224_ ) );
OAI21_X1 \RegFile/_7756_ ( .A(\RegFile/_3224_ ), .B1(\RegFile/_2399_ ), .B2(\RegFile/_3209_ ), .ZN(\RegFile/_0558_ ) );
AOI21_X1 \RegFile/_7757_ ( .A(\RegFile/_2404_ ), .B1(\RegFile/_2417_ ), .B2(\RegFile/_2418_ ), .ZN(\RegFile/_3225_ ) );
AOI21_X1 \RegFile/_7758_ ( .A(\RegFile/_3225_ ), .B1(\RegFile/_1097_ ), .B2(\RegFile/_3209_ ), .ZN(\RegFile/_0559_ ) );
NAND3_X1 \RegFile/_7759_ ( .A1(\RegFile/_2437_ ), .A2(\RegFile/_2031_ ), .A3(\RegFile/_2438_ ), .ZN(\RegFile/_3226_ ) );
BUF_X4 \RegFile/_7760_ ( .A(\RegFile/_2031_ ), .Z(\RegFile/_3227_ ) );
OAI21_X1 \RegFile/_7761_ ( .A(\RegFile/_3226_ ), .B1(\RegFile/_1734_ ), .B2(\RegFile/_3227_ ), .ZN(\RegFile/_0560_ ) );
NAND2_X1 \RegFile/_7762_ ( .A1(\RegFile/_3212_ ), .A2(\RegFile/_3418_ ), .ZN(\RegFile/_3228_ ) );
OAI21_X1 \RegFile/_7763_ ( .A(\RegFile/_3228_ ), .B1(\RegFile/_2458_ ), .B2(\RegFile/_3209_ ), .ZN(\RegFile/_0561_ ) );
NAND2_X1 \RegFile/_7764_ ( .A1(\RegFile/_3212_ ), .A2(\RegFile/_3419_ ), .ZN(\RegFile/_3229_ ) );
OAI21_X1 \RegFile/_7765_ ( .A(\RegFile/_3229_ ), .B1(\RegFile/_2476_ ), .B2(\RegFile/_3209_ ), .ZN(\RegFile/_0562_ ) );
OR3_X1 \RegFile/_7766_ ( .A1(\RegFile/_2492_ ), .A2(\RegFile/_2404_ ), .A3(\RegFile/_2493_ ), .ZN(\RegFile/_3230_ ) );
OAI21_X1 \RegFile/_7767_ ( .A(\RegFile/_3230_ ), .B1(\RegFile/_1164_ ), .B2(\RegFile/_3227_ ), .ZN(\RegFile/_0563_ ) );
OR3_X1 \RegFile/_7768_ ( .A1(\RegFile/_2511_ ), .A2(\RegFile/_2404_ ), .A3(\RegFile/_2512_ ), .ZN(\RegFile/_3231_ ) );
OAI21_X1 \RegFile/_7769_ ( .A(\RegFile/_3231_ ), .B1(\RegFile/_1184_ ), .B2(\RegFile/_3227_ ), .ZN(\RegFile/_0564_ ) );
AOI21_X1 \RegFile/_7770_ ( .A(\RegFile/_3423_ ), .B1(\RegFile/_3210_ ), .B2(\RegFile/_3165_ ), .ZN(\RegFile/_3232_ ) );
AOI21_X1 \RegFile/_7771_ ( .A(\RegFile/_3232_ ), .B1(\RegFile/_2533_ ), .B2(\RegFile/_3207_ ), .ZN(\RegFile/_0565_ ) );
NAND2_X1 \RegFile/_7772_ ( .A1(\RegFile/_3212_ ), .A2(\RegFile/_3424_ ), .ZN(\RegFile/_3233_ ) );
OAI21_X1 \RegFile/_7773_ ( .A(\RegFile/_3233_ ), .B1(\RegFile/_2551_ ), .B2(\RegFile/_3209_ ), .ZN(\RegFile/_0566_ ) );
NAND2_X1 \RegFile/_7774_ ( .A1(\RegFile/_2404_ ), .A2(\RegFile/_3425_ ), .ZN(\RegFile/_3234_ ) );
OAI21_X1 \RegFile/_7775_ ( .A(\RegFile/_3234_ ), .B1(\RegFile/_2570_ ), .B2(\RegFile/_3212_ ), .ZN(\RegFile/_0567_ ) );
NAND3_X1 \RegFile/_7776_ ( .A1(\RegFile/_2589_ ), .A2(\RegFile/_2031_ ), .A3(\RegFile/_2590_ ), .ZN(\RegFile/_3235_ ) );
OAI21_X1 \RegFile/_7777_ ( .A(\RegFile/_3235_ ), .B1(\RegFile/_1249_ ), .B2(\RegFile/_3227_ ), .ZN(\RegFile/_0568_ ) );
AOI21_X1 \RegFile/_7778_ ( .A(\RegFile/_3427_ ), .B1(\RegFile/_3210_ ), .B2(\RegFile/_3165_ ), .ZN(\RegFile/_3236_ ) );
AOI21_X1 \RegFile/_7779_ ( .A(\RegFile/_3236_ ), .B1(\RegFile/_2608_ ), .B2(\RegFile/_3227_ ), .ZN(\RegFile/_0569_ ) );
AOI21_X1 \RegFile/_7780_ ( .A(\RegFile/_3428_ ), .B1(\RegFile/_3045_ ), .B2(\RegFile/_3165_ ), .ZN(\RegFile/_3237_ ) );
AOI21_X1 \RegFile/_7781_ ( .A(\RegFile/_3237_ ), .B1(\RegFile/_2628_ ), .B2(\RegFile/_3227_ ), .ZN(\RegFile/_0570_ ) );
AOI21_X1 \RegFile/_7782_ ( .A(\RegFile/_3429_ ), .B1(\RegFile/_3045_ ), .B2(\RegFile/_3165_ ), .ZN(\RegFile/_3238_ ) );
AOI21_X1 \RegFile/_7783_ ( .A(\RegFile/_3238_ ), .B1(\RegFile/_2646_ ), .B2(\RegFile/_3227_ ), .ZN(\RegFile/_0571_ ) );
AOI21_X1 \RegFile/_7784_ ( .A(\RegFile/_3430_ ), .B1(\RegFile/_3045_ ), .B2(\RegFile/_3165_ ), .ZN(\RegFile/_3239_ ) );
AOI21_X1 \RegFile/_7785_ ( .A(\RegFile/_3239_ ), .B1(\RegFile/_2664_ ), .B2(\RegFile/_3227_ ), .ZN(\RegFile/_0572_ ) );
AOI21_X1 \RegFile/_7786_ ( .A(\RegFile/_3431_ ), .B1(\RegFile/_3045_ ), .B2(\RegFile/_3165_ ), .ZN(\RegFile/_3240_ ) );
AOI21_X1 \RegFile/_7787_ ( .A(\RegFile/_3240_ ), .B1(\RegFile/_2685_ ), .B2(\RegFile/_3227_ ), .ZN(\RegFile/_0573_ ) );
NAND2_X1 \RegFile/_7788_ ( .A1(\RegFile/_2404_ ), .A2(\RegFile/_3433_ ), .ZN(\RegFile/_3241_ ) );
OAI21_X1 \RegFile/_7789_ ( .A(\RegFile/_3241_ ), .B1(\RegFile/_2704_ ), .B2(\RegFile/_3212_ ), .ZN(\RegFile/_0574_ ) );
AOI21_X1 \RegFile/_7790_ ( .A(\RegFile/_3434_ ), .B1(\RegFile/_3045_ ), .B2(\RegFile/_3165_ ), .ZN(\RegFile/_3242_ ) );
AOI21_X1 \RegFile/_7791_ ( .A(\RegFile/_3242_ ), .B1(\RegFile/_2723_ ), .B2(\RegFile/_3227_ ), .ZN(\RegFile/_0575_ ) );
NAND2_X2 \RegFile/_7792_ ( .A1(\RegFile/_2169_ ), .A2(\RegFile/_1996_ ), .ZN(\RegFile/_3243_ ) );
BUF_X4 \RegFile/_7793_ ( .A(\RegFile/_3243_ ), .Z(\RegFile/_3244_ ) );
NAND2_X1 \RegFile/_7794_ ( .A1(\RegFile/_3244_ ), .A2(\RegFile/_3442_ ), .ZN(\RegFile/_3245_ ) );
BUF_X4 \RegFile/_7795_ ( .A(\RegFile/_3243_ ), .Z(\RegFile/_3246_ ) );
OAI21_X1 \RegFile/_7796_ ( .A(\RegFile/_3245_ ), .B1(\RegFile/_2071_ ), .B2(\RegFile/_3246_ ), .ZN(\RegFile/_0576_ ) );
NAND2_X1 \RegFile/_7797_ ( .A1(\RegFile/_3244_ ), .A2(\RegFile/_3453_ ), .ZN(\RegFile/_3247_ ) );
OAI21_X1 \RegFile/_7798_ ( .A(\RegFile/_3247_ ), .B1(\RegFile/_2112_ ), .B2(\RegFile/_3246_ ), .ZN(\RegFile/_0577_ ) );
NAND2_X1 \RegFile/_7799_ ( .A1(\RegFile/_3244_ ), .A2(\RegFile/_3464_ ), .ZN(\RegFile/_3248_ ) );
OAI21_X1 \RegFile/_7800_ ( .A(\RegFile/_3248_ ), .B1(\RegFile/_2141_ ), .B2(\RegFile/_3246_ ), .ZN(\RegFile/_0578_ ) );
NAND2_X1 \RegFile/_7801_ ( .A1(\RegFile/_3244_ ), .A2(\RegFile/_3467_ ), .ZN(\RegFile/_3249_ ) );
OAI21_X1 \RegFile/_7802_ ( .A(\RegFile/_3249_ ), .B1(\RegFile/_2175_ ), .B2(\RegFile/_3246_ ), .ZN(\RegFile/_0579_ ) );
NAND2_X1 \RegFile/_7803_ ( .A1(\RegFile/_3244_ ), .A2(\RegFile/_3468_ ), .ZN(\RegFile/_3250_ ) );
OAI21_X1 \RegFile/_7804_ ( .A(\RegFile/_3250_ ), .B1(\RegFile/_2198_ ), .B2(\RegFile/_3246_ ), .ZN(\RegFile/_0580_ ) );
NAND2_X1 \RegFile/_7805_ ( .A1(\RegFile/_3244_ ), .A2(\RegFile/_3469_ ), .ZN(\RegFile/_3251_ ) );
OAI21_X1 \RegFile/_7806_ ( .A(\RegFile/_3251_ ), .B1(\RegFile/_2218_ ), .B2(\RegFile/_3246_ ), .ZN(\RegFile/_0581_ ) );
NAND2_X1 \RegFile/_7807_ ( .A1(\RegFile/_3244_ ), .A2(\RegFile/_3470_ ), .ZN(\RegFile/_3252_ ) );
OAI21_X1 \RegFile/_7808_ ( .A(\RegFile/_3252_ ), .B1(\RegFile/_2239_ ), .B2(\RegFile/_3246_ ), .ZN(\RegFile/_0582_ ) );
NAND2_X1 \RegFile/_7809_ ( .A1(\RegFile/_3244_ ), .A2(\RegFile/_3471_ ), .ZN(\RegFile/_3253_ ) );
OAI21_X1 \RegFile/_7810_ ( .A(\RegFile/_3253_ ), .B1(\RegFile/_2260_ ), .B2(\RegFile/_3246_ ), .ZN(\RegFile/_0583_ ) );
BUF_X4 \RegFile/_7811_ ( .A(\RegFile/_3243_ ), .Z(\RegFile/_3254_ ) );
NAND2_X1 \RegFile/_7812_ ( .A1(\RegFile/_3254_ ), .A2(\RegFile/_3472_ ), .ZN(\RegFile/_3255_ ) );
OAI21_X1 \RegFile/_7813_ ( .A(\RegFile/_3255_ ), .B1(\RegFile/_2280_ ), .B2(\RegFile/_3246_ ), .ZN(\RegFile/_0584_ ) );
NAND2_X1 \RegFile/_7814_ ( .A1(\RegFile/_3254_ ), .A2(\RegFile/_3473_ ), .ZN(\RegFile/_3256_ ) );
OAI21_X1 \RegFile/_7815_ ( .A(\RegFile/_3256_ ), .B1(\RegFile/_2298_ ), .B2(\RegFile/_3246_ ), .ZN(\RegFile/_0585_ ) );
NAND2_X1 \RegFile/_7816_ ( .A1(\RegFile/_3254_ ), .A2(\RegFile/_3443_ ), .ZN(\RegFile/_3257_ ) );
BUF_X4 \RegFile/_7817_ ( .A(\RegFile/_3243_ ), .Z(\RegFile/_3258_ ) );
OAI21_X1 \RegFile/_7818_ ( .A(\RegFile/_3257_ ), .B1(\RegFile/_2317_ ), .B2(\RegFile/_3258_ ), .ZN(\RegFile/_0586_ ) );
NAND2_X1 \RegFile/_7819_ ( .A1(\RegFile/_3254_ ), .A2(\RegFile/_3444_ ), .ZN(\RegFile/_3259_ ) );
OAI21_X1 \RegFile/_7820_ ( .A(\RegFile/_3259_ ), .B1(\RegFile/_2335_ ), .B2(\RegFile/_3258_ ), .ZN(\RegFile/_0587_ ) );
NAND2_X1 \RegFile/_7821_ ( .A1(\RegFile/_3254_ ), .A2(\RegFile/_3445_ ), .ZN(\RegFile/_3260_ ) );
OAI21_X1 \RegFile/_7822_ ( .A(\RegFile/_3260_ ), .B1(\RegFile/_2356_ ), .B2(\RegFile/_3258_ ), .ZN(\RegFile/_0588_ ) );
NAND2_X1 \RegFile/_7823_ ( .A1(\RegFile/_3254_ ), .A2(\RegFile/_3446_ ), .ZN(\RegFile/_3261_ ) );
OAI21_X1 \RegFile/_7824_ ( .A(\RegFile/_3261_ ), .B1(\RegFile/_2378_ ), .B2(\RegFile/_3258_ ), .ZN(\RegFile/_0589_ ) );
NAND2_X1 \RegFile/_7825_ ( .A1(\RegFile/_3254_ ), .A2(\RegFile/_3447_ ), .ZN(\RegFile/_3262_ ) );
OAI21_X1 \RegFile/_7826_ ( .A(\RegFile/_3262_ ), .B1(\RegFile/_2399_ ), .B2(\RegFile/_3258_ ), .ZN(\RegFile/_0590_ ) );
NAND2_X1 \RegFile/_7827_ ( .A1(\RegFile/_3254_ ), .A2(\RegFile/_3448_ ), .ZN(\RegFile/_3263_ ) );
OAI21_X1 \RegFile/_7828_ ( .A(\RegFile/_3263_ ), .B1(\RegFile/_2419_ ), .B2(\RegFile/_3258_ ), .ZN(\RegFile/_0591_ ) );
NAND2_X1 \RegFile/_7829_ ( .A1(\RegFile/_3254_ ), .A2(\RegFile/_3449_ ), .ZN(\RegFile/_3264_ ) );
OAI21_X1 \RegFile/_7830_ ( .A(\RegFile/_3264_ ), .B1(\RegFile/_2439_ ), .B2(\RegFile/_3258_ ), .ZN(\RegFile/_0592_ ) );
NAND2_X1 \RegFile/_7831_ ( .A1(\RegFile/_3254_ ), .A2(\RegFile/_3450_ ), .ZN(\RegFile/_3265_ ) );
OAI21_X1 \RegFile/_7832_ ( .A(\RegFile/_3265_ ), .B1(\RegFile/_2458_ ), .B2(\RegFile/_3258_ ), .ZN(\RegFile/_0593_ ) );
BUF_X4 \RegFile/_7833_ ( .A(\RegFile/_3243_ ), .Z(\RegFile/_3266_ ) );
NAND2_X1 \RegFile/_7834_ ( .A1(\RegFile/_3266_ ), .A2(\RegFile/_3451_ ), .ZN(\RegFile/_3267_ ) );
OAI21_X1 \RegFile/_7835_ ( .A(\RegFile/_3267_ ), .B1(\RegFile/_2475_ ), .B2(\RegFile/_3258_ ), .ZN(\RegFile/_0594_ ) );
NAND2_X1 \RegFile/_7836_ ( .A1(\RegFile/_3266_ ), .A2(\RegFile/_3452_ ), .ZN(\RegFile/_3268_ ) );
OAI21_X1 \RegFile/_7837_ ( .A(\RegFile/_3268_ ), .B1(\RegFile/_2495_ ), .B2(\RegFile/_3258_ ), .ZN(\RegFile/_0595_ ) );
NAND2_X1 \RegFile/_7838_ ( .A1(\RegFile/_3266_ ), .A2(\RegFile/_3454_ ), .ZN(\RegFile/_3269_ ) );
BUF_X4 \RegFile/_7839_ ( .A(\RegFile/_3243_ ), .Z(\RegFile/_3270_ ) );
OAI21_X1 \RegFile/_7840_ ( .A(\RegFile/_3269_ ), .B1(\RegFile/_2514_ ), .B2(\RegFile/_3270_ ), .ZN(\RegFile/_0596_ ) );
NAND2_X1 \RegFile/_7841_ ( .A1(\RegFile/_3266_ ), .A2(\RegFile/_3455_ ), .ZN(\RegFile/_3271_ ) );
OAI21_X1 \RegFile/_7842_ ( .A(\RegFile/_3271_ ), .B1(\RegFile/_2532_ ), .B2(\RegFile/_3270_ ), .ZN(\RegFile/_0597_ ) );
NAND2_X1 \RegFile/_7843_ ( .A1(\RegFile/_3266_ ), .A2(\RegFile/_3456_ ), .ZN(\RegFile/_3272_ ) );
OAI21_X1 \RegFile/_7844_ ( .A(\RegFile/_3272_ ), .B1(\RegFile/_2551_ ), .B2(\RegFile/_3270_ ), .ZN(\RegFile/_0598_ ) );
NAND2_X1 \RegFile/_7845_ ( .A1(\RegFile/_3266_ ), .A2(\RegFile/_3457_ ), .ZN(\RegFile/_3273_ ) );
OAI21_X1 \RegFile/_7846_ ( .A(\RegFile/_3273_ ), .B1(\RegFile/_2570_ ), .B2(\RegFile/_3270_ ), .ZN(\RegFile/_0599_ ) );
NAND2_X1 \RegFile/_7847_ ( .A1(\RegFile/_3266_ ), .A2(\RegFile/_3458_ ), .ZN(\RegFile/_3274_ ) );
OAI21_X1 \RegFile/_7848_ ( .A(\RegFile/_3274_ ), .B1(\RegFile/_2591_ ), .B2(\RegFile/_3270_ ), .ZN(\RegFile/_0600_ ) );
NAND2_X1 \RegFile/_7849_ ( .A1(\RegFile/_3266_ ), .A2(\RegFile/_3459_ ), .ZN(\RegFile/_3275_ ) );
OAI21_X1 \RegFile/_7850_ ( .A(\RegFile/_3275_ ), .B1(\RegFile/_2608_ ), .B2(\RegFile/_3270_ ), .ZN(\RegFile/_0601_ ) );
NAND2_X1 \RegFile/_7851_ ( .A1(\RegFile/_3266_ ), .A2(\RegFile/_3460_ ), .ZN(\RegFile/_3276_ ) );
OAI21_X1 \RegFile/_7852_ ( .A(\RegFile/_3276_ ), .B1(\RegFile/_2627_ ), .B2(\RegFile/_3270_ ), .ZN(\RegFile/_0602_ ) );
NAND2_X1 \RegFile/_7853_ ( .A1(\RegFile/_3266_ ), .A2(\RegFile/_3461_ ), .ZN(\RegFile/_3277_ ) );
OAI21_X1 \RegFile/_7854_ ( .A(\RegFile/_3277_ ), .B1(\RegFile/_2645_ ), .B2(\RegFile/_3270_ ), .ZN(\RegFile/_0603_ ) );
NAND2_X1 \RegFile/_7855_ ( .A1(\RegFile/_3243_ ), .A2(\RegFile/_3462_ ), .ZN(\RegFile/_3278_ ) );
OAI21_X1 \RegFile/_7856_ ( .A(\RegFile/_3278_ ), .B1(\RegFile/_2663_ ), .B2(\RegFile/_3270_ ), .ZN(\RegFile/_0604_ ) );
NAND2_X1 \RegFile/_7857_ ( .A1(\RegFile/_3243_ ), .A2(\RegFile/_3463_ ), .ZN(\RegFile/_3279_ ) );
OAI21_X1 \RegFile/_7858_ ( .A(\RegFile/_3279_ ), .B1(\RegFile/_2684_ ), .B2(\RegFile/_3270_ ), .ZN(\RegFile/_0605_ ) );
NAND2_X1 \RegFile/_7859_ ( .A1(\RegFile/_3243_ ), .A2(\RegFile/_3465_ ), .ZN(\RegFile/_3280_ ) );
OAI21_X1 \RegFile/_7860_ ( .A(\RegFile/_3280_ ), .B1(\RegFile/_2704_ ), .B2(\RegFile/_3244_ ), .ZN(\RegFile/_0606_ ) );
NAND2_X1 \RegFile/_7861_ ( .A1(\RegFile/_3243_ ), .A2(\RegFile/_3466_ ), .ZN(\RegFile/_3281_ ) );
OAI21_X1 \RegFile/_7862_ ( .A(\RegFile/_3281_ ), .B1(\RegFile/_2723_ ), .B2(\RegFile/_3244_ ), .ZN(\RegFile/_0607_ ) );
DFF_X1 \RegFile/_7863_ ( .D(\RegFile/_4242_ ), .CK(clock ), .Q(\RegFile/reg_0 [0] ), .QN(\RegFile/_4241_ ) );
DFF_X1 \RegFile/_7864_ ( .D(\RegFile/_4243_ ), .CK(clock ), .Q(\RegFile/reg_0 [1] ), .QN(\RegFile/_4240_ ) );
DFF_X1 \RegFile/_7865_ ( .D(\RegFile/_4244_ ), .CK(clock ), .Q(\RegFile/reg_0 [2] ), .QN(\RegFile/_4239_ ) );
DFF_X1 \RegFile/_7866_ ( .D(\RegFile/_4245_ ), .CK(clock ), .Q(\RegFile/reg_0 [3] ), .QN(\RegFile/_4238_ ) );
DFF_X1 \RegFile/_7867_ ( .D(\RegFile/_4246_ ), .CK(clock ), .Q(\RegFile/reg_0 [4] ), .QN(\RegFile/_4237_ ) );
DFF_X1 \RegFile/_7868_ ( .D(\RegFile/_4247_ ), .CK(clock ), .Q(\RegFile/reg_0 [5] ), .QN(\RegFile/_4236_ ) );
DFF_X1 \RegFile/_7869_ ( .D(\RegFile/_4248_ ), .CK(clock ), .Q(\RegFile/reg_0 [6] ), .QN(\RegFile/_4235_ ) );
DFF_X1 \RegFile/_7870_ ( .D(\RegFile/_4249_ ), .CK(clock ), .Q(\RegFile/reg_0 [7] ), .QN(\RegFile/_4234_ ) );
DFF_X1 \RegFile/_7871_ ( .D(\RegFile/_4250_ ), .CK(clock ), .Q(\RegFile/reg_0 [8] ), .QN(\RegFile/_4233_ ) );
DFF_X1 \RegFile/_7872_ ( .D(\RegFile/_4251_ ), .CK(clock ), .Q(\RegFile/reg_0 [9] ), .QN(\RegFile/_4232_ ) );
DFF_X1 \RegFile/_7873_ ( .D(\RegFile/_4252_ ), .CK(clock ), .Q(\RegFile/reg_0 [10] ), .QN(\RegFile/_4231_ ) );
DFF_X1 \RegFile/_7874_ ( .D(\RegFile/_4253_ ), .CK(clock ), .Q(\RegFile/reg_0 [11] ), .QN(\RegFile/_4230_ ) );
DFF_X1 \RegFile/_7875_ ( .D(\RegFile/_4254_ ), .CK(clock ), .Q(\RegFile/reg_0 [12] ), .QN(\RegFile/_4229_ ) );
DFF_X1 \RegFile/_7876_ ( .D(\RegFile/_4255_ ), .CK(clock ), .Q(\RegFile/reg_0 [13] ), .QN(\RegFile/_4228_ ) );
DFF_X1 \RegFile/_7877_ ( .D(\RegFile/_4256_ ), .CK(clock ), .Q(\RegFile/reg_0 [14] ), .QN(\RegFile/_4227_ ) );
DFF_X1 \RegFile/_7878_ ( .D(\RegFile/_4257_ ), .CK(clock ), .Q(\RegFile/reg_0 [15] ), .QN(\RegFile/_4226_ ) );
DFF_X1 \RegFile/_7879_ ( .D(\RegFile/_4258_ ), .CK(clock ), .Q(\RegFile/reg_0 [16] ), .QN(\RegFile/_4225_ ) );
DFF_X1 \RegFile/_7880_ ( .D(\RegFile/_4259_ ), .CK(clock ), .Q(\RegFile/reg_0 [17] ), .QN(\RegFile/_4224_ ) );
DFF_X1 \RegFile/_7881_ ( .D(\RegFile/_4260_ ), .CK(clock ), .Q(\RegFile/reg_0 [18] ), .QN(\RegFile/_4223_ ) );
DFF_X1 \RegFile/_7882_ ( .D(\RegFile/_4261_ ), .CK(clock ), .Q(\RegFile/reg_0 [19] ), .QN(\RegFile/_4222_ ) );
DFF_X1 \RegFile/_7883_ ( .D(\RegFile/_4262_ ), .CK(clock ), .Q(\RegFile/reg_0 [20] ), .QN(\RegFile/_4221_ ) );
DFF_X1 \RegFile/_7884_ ( .D(\RegFile/_4263_ ), .CK(clock ), .Q(\RegFile/reg_0 [21] ), .QN(\RegFile/_4220_ ) );
DFF_X1 \RegFile/_7885_ ( .D(\RegFile/_4264_ ), .CK(clock ), .Q(\RegFile/reg_0 [22] ), .QN(\RegFile/_4219_ ) );
DFF_X1 \RegFile/_7886_ ( .D(\RegFile/_4265_ ), .CK(clock ), .Q(\RegFile/reg_0 [23] ), .QN(\RegFile/_4218_ ) );
DFF_X1 \RegFile/_7887_ ( .D(\RegFile/_4266_ ), .CK(clock ), .Q(\RegFile/reg_0 [24] ), .QN(\RegFile/_4217_ ) );
DFF_X1 \RegFile/_7888_ ( .D(\RegFile/_4267_ ), .CK(clock ), .Q(\RegFile/reg_0 [25] ), .QN(\RegFile/_4216_ ) );
DFF_X1 \RegFile/_7889_ ( .D(\RegFile/_4268_ ), .CK(clock ), .Q(\RegFile/reg_0 [26] ), .QN(\RegFile/_4215_ ) );
DFF_X1 \RegFile/_7890_ ( .D(\RegFile/_4269_ ), .CK(clock ), .Q(\RegFile/reg_0 [27] ), .QN(\RegFile/_4214_ ) );
DFF_X1 \RegFile/_7891_ ( .D(\RegFile/_4270_ ), .CK(clock ), .Q(\RegFile/reg_0 [28] ), .QN(\RegFile/_4213_ ) );
DFF_X1 \RegFile/_7892_ ( .D(\RegFile/_4271_ ), .CK(clock ), .Q(\RegFile/reg_0 [29] ), .QN(\RegFile/_4212_ ) );
DFF_X1 \RegFile/_7893_ ( .D(\RegFile/_4272_ ), .CK(clock ), .Q(\RegFile/reg_0 [30] ), .QN(\RegFile/_4211_ ) );
DFF_X1 \RegFile/_7894_ ( .D(\RegFile/_4273_ ), .CK(clock ), .Q(\RegFile/reg_0 [31] ), .QN(\RegFile/_4210_ ) );
DFF_X1 \RegFile/_7895_ ( .D(\RegFile/_4274_ ), .CK(clock ), .Q(\RegFile/reg_1 [0] ), .QN(\RegFile/_4209_ ) );
DFF_X1 \RegFile/_7896_ ( .D(\RegFile/_4275_ ), .CK(clock ), .Q(\RegFile/reg_1 [1] ), .QN(\RegFile/_4208_ ) );
DFF_X1 \RegFile/_7897_ ( .D(\RegFile/_4276_ ), .CK(clock ), .Q(\RegFile/reg_1 [2] ), .QN(\RegFile/_4207_ ) );
DFF_X1 \RegFile/_7898_ ( .D(\RegFile/_4277_ ), .CK(clock ), .Q(\RegFile/reg_1 [3] ), .QN(\RegFile/_4206_ ) );
DFF_X1 \RegFile/_7899_ ( .D(\RegFile/_4278_ ), .CK(clock ), .Q(\RegFile/reg_1 [4] ), .QN(\RegFile/_4205_ ) );
DFF_X1 \RegFile/_7900_ ( .D(\RegFile/_4279_ ), .CK(clock ), .Q(\RegFile/reg_1 [5] ), .QN(\RegFile/_4204_ ) );
DFF_X1 \RegFile/_7901_ ( .D(\RegFile/_4280_ ), .CK(clock ), .Q(\RegFile/reg_1 [6] ), .QN(\RegFile/_4203_ ) );
DFF_X1 \RegFile/_7902_ ( .D(\RegFile/_4281_ ), .CK(clock ), .Q(\RegFile/reg_1 [7] ), .QN(\RegFile/_4202_ ) );
DFF_X1 \RegFile/_7903_ ( .D(\RegFile/_4282_ ), .CK(clock ), .Q(\RegFile/reg_1 [8] ), .QN(\RegFile/_4201_ ) );
DFF_X1 \RegFile/_7904_ ( .D(\RegFile/_4283_ ), .CK(clock ), .Q(\RegFile/reg_1 [9] ), .QN(\RegFile/_4200_ ) );
DFF_X1 \RegFile/_7905_ ( .D(\RegFile/_4284_ ), .CK(clock ), .Q(\RegFile/reg_1 [10] ), .QN(\RegFile/_4199_ ) );
DFF_X1 \RegFile/_7906_ ( .D(\RegFile/_4285_ ), .CK(clock ), .Q(\RegFile/reg_1 [11] ), .QN(\RegFile/_4198_ ) );
DFF_X1 \RegFile/_7907_ ( .D(\RegFile/_4286_ ), .CK(clock ), .Q(\RegFile/reg_1 [12] ), .QN(\RegFile/_4197_ ) );
DFF_X1 \RegFile/_7908_ ( .D(\RegFile/_4287_ ), .CK(clock ), .Q(\RegFile/reg_1 [13] ), .QN(\RegFile/_4196_ ) );
DFF_X1 \RegFile/_7909_ ( .D(\RegFile/_4288_ ), .CK(clock ), .Q(\RegFile/reg_1 [14] ), .QN(\RegFile/_4195_ ) );
DFF_X1 \RegFile/_7910_ ( .D(\RegFile/_4289_ ), .CK(clock ), .Q(\RegFile/reg_1 [15] ), .QN(\RegFile/_4194_ ) );
DFF_X1 \RegFile/_7911_ ( .D(\RegFile/_4290_ ), .CK(clock ), .Q(\RegFile/reg_1 [16] ), .QN(\RegFile/_4193_ ) );
DFF_X1 \RegFile/_7912_ ( .D(\RegFile/_4291_ ), .CK(clock ), .Q(\RegFile/reg_1 [17] ), .QN(\RegFile/_4192_ ) );
DFF_X1 \RegFile/_7913_ ( .D(\RegFile/_4292_ ), .CK(clock ), .Q(\RegFile/reg_1 [18] ), .QN(\RegFile/_4191_ ) );
DFF_X1 \RegFile/_7914_ ( .D(\RegFile/_4293_ ), .CK(clock ), .Q(\RegFile/reg_1 [19] ), .QN(\RegFile/_4190_ ) );
DFF_X1 \RegFile/_7915_ ( .D(\RegFile/_4294_ ), .CK(clock ), .Q(\RegFile/reg_1 [20] ), .QN(\RegFile/_4189_ ) );
DFF_X1 \RegFile/_7916_ ( .D(\RegFile/_4295_ ), .CK(clock ), .Q(\RegFile/reg_1 [21] ), .QN(\RegFile/_4188_ ) );
DFF_X1 \RegFile/_7917_ ( .D(\RegFile/_4296_ ), .CK(clock ), .Q(\RegFile/reg_1 [22] ), .QN(\RegFile/_4187_ ) );
DFF_X1 \RegFile/_7918_ ( .D(\RegFile/_4297_ ), .CK(clock ), .Q(\RegFile/reg_1 [23] ), .QN(\RegFile/_4186_ ) );
DFF_X1 \RegFile/_7919_ ( .D(\RegFile/_4298_ ), .CK(clock ), .Q(\RegFile/reg_1 [24] ), .QN(\RegFile/_4185_ ) );
DFF_X1 \RegFile/_7920_ ( .D(\RegFile/_4299_ ), .CK(clock ), .Q(\RegFile/reg_1 [25] ), .QN(\RegFile/_4184_ ) );
DFF_X1 \RegFile/_7921_ ( .D(\RegFile/_4300_ ), .CK(clock ), .Q(\RegFile/reg_1 [26] ), .QN(\RegFile/_4183_ ) );
DFF_X1 \RegFile/_7922_ ( .D(\RegFile/_4301_ ), .CK(clock ), .Q(\RegFile/reg_1 [27] ), .QN(\RegFile/_4182_ ) );
DFF_X1 \RegFile/_7923_ ( .D(\RegFile/_4302_ ), .CK(clock ), .Q(\RegFile/reg_1 [28] ), .QN(\RegFile/_4181_ ) );
DFF_X1 \RegFile/_7924_ ( .D(\RegFile/_4303_ ), .CK(clock ), .Q(\RegFile/reg_1 [29] ), .QN(\RegFile/_4180_ ) );
DFF_X1 \RegFile/_7925_ ( .D(\RegFile/_4304_ ), .CK(clock ), .Q(\RegFile/reg_1 [30] ), .QN(\RegFile/_4179_ ) );
DFF_X1 \RegFile/_7926_ ( .D(\RegFile/_4305_ ), .CK(clock ), .Q(\RegFile/reg_1 [31] ), .QN(\RegFile/_4178_ ) );
DFF_X1 \RegFile/_7927_ ( .D(\RegFile/_4306_ ), .CK(clock ), .Q(\RegFile/reg_2 [0] ), .QN(\RegFile/_4177_ ) );
DFF_X1 \RegFile/_7928_ ( .D(\RegFile/_4307_ ), .CK(clock ), .Q(\RegFile/reg_2 [1] ), .QN(\RegFile/_4176_ ) );
DFF_X1 \RegFile/_7929_ ( .D(\RegFile/_4308_ ), .CK(clock ), .Q(\RegFile/reg_2 [2] ), .QN(\RegFile/_4175_ ) );
DFF_X1 \RegFile/_7930_ ( .D(\RegFile/_4309_ ), .CK(clock ), .Q(\RegFile/reg_2 [3] ), .QN(\RegFile/_4174_ ) );
DFF_X1 \RegFile/_7931_ ( .D(\RegFile/_4310_ ), .CK(clock ), .Q(\RegFile/reg_2 [4] ), .QN(\RegFile/_4173_ ) );
DFF_X1 \RegFile/_7932_ ( .D(\RegFile/_4311_ ), .CK(clock ), .Q(\RegFile/reg_2 [5] ), .QN(\RegFile/_4172_ ) );
DFF_X1 \RegFile/_7933_ ( .D(\RegFile/_4312_ ), .CK(clock ), .Q(\RegFile/reg_2 [6] ), .QN(\RegFile/_4171_ ) );
DFF_X1 \RegFile/_7934_ ( .D(\RegFile/_4313_ ), .CK(clock ), .Q(\RegFile/reg_2 [7] ), .QN(\RegFile/_4170_ ) );
DFF_X1 \RegFile/_7935_ ( .D(\RegFile/_4314_ ), .CK(clock ), .Q(\RegFile/reg_2 [8] ), .QN(\RegFile/_4169_ ) );
DFF_X1 \RegFile/_7936_ ( .D(\RegFile/_4315_ ), .CK(clock ), .Q(\RegFile/reg_2 [9] ), .QN(\RegFile/_4168_ ) );
DFF_X1 \RegFile/_7937_ ( .D(\RegFile/_4316_ ), .CK(clock ), .Q(\RegFile/reg_2 [10] ), .QN(\RegFile/_4167_ ) );
DFF_X1 \RegFile/_7938_ ( .D(\RegFile/_4317_ ), .CK(clock ), .Q(\RegFile/reg_2 [11] ), .QN(\RegFile/_4166_ ) );
DFF_X1 \RegFile/_7939_ ( .D(\RegFile/_4318_ ), .CK(clock ), .Q(\RegFile/reg_2 [12] ), .QN(\RegFile/_4165_ ) );
DFF_X1 \RegFile/_7940_ ( .D(\RegFile/_4319_ ), .CK(clock ), .Q(\RegFile/reg_2 [13] ), .QN(\RegFile/_4164_ ) );
DFF_X1 \RegFile/_7941_ ( .D(\RegFile/_4320_ ), .CK(clock ), .Q(\RegFile/reg_2 [14] ), .QN(\RegFile/_4163_ ) );
DFF_X1 \RegFile/_7942_ ( .D(\RegFile/_4321_ ), .CK(clock ), .Q(\RegFile/reg_2 [15] ), .QN(\RegFile/_4162_ ) );
DFF_X1 \RegFile/_7943_ ( .D(\RegFile/_4322_ ), .CK(clock ), .Q(\RegFile/reg_2 [16] ), .QN(\RegFile/_4161_ ) );
DFF_X1 \RegFile/_7944_ ( .D(\RegFile/_4323_ ), .CK(clock ), .Q(\RegFile/reg_2 [17] ), .QN(\RegFile/_4160_ ) );
DFF_X1 \RegFile/_7945_ ( .D(\RegFile/_4324_ ), .CK(clock ), .Q(\RegFile/reg_2 [18] ), .QN(\RegFile/_4159_ ) );
DFF_X1 \RegFile/_7946_ ( .D(\RegFile/_4325_ ), .CK(clock ), .Q(\RegFile/reg_2 [19] ), .QN(\RegFile/_4158_ ) );
DFF_X1 \RegFile/_7947_ ( .D(\RegFile/_4326_ ), .CK(clock ), .Q(\RegFile/reg_2 [20] ), .QN(\RegFile/_4157_ ) );
DFF_X1 \RegFile/_7948_ ( .D(\RegFile/_4327_ ), .CK(clock ), .Q(\RegFile/reg_2 [21] ), .QN(\RegFile/_4156_ ) );
DFF_X1 \RegFile/_7949_ ( .D(\RegFile/_4328_ ), .CK(clock ), .Q(\RegFile/reg_2 [22] ), .QN(\RegFile/_4155_ ) );
DFF_X1 \RegFile/_7950_ ( .D(\RegFile/_4329_ ), .CK(clock ), .Q(\RegFile/reg_2 [23] ), .QN(\RegFile/_4154_ ) );
DFF_X1 \RegFile/_7951_ ( .D(\RegFile/_4330_ ), .CK(clock ), .Q(\RegFile/reg_2 [24] ), .QN(\RegFile/_4153_ ) );
DFF_X1 \RegFile/_7952_ ( .D(\RegFile/_4331_ ), .CK(clock ), .Q(\RegFile/reg_2 [25] ), .QN(\RegFile/_4152_ ) );
DFF_X1 \RegFile/_7953_ ( .D(\RegFile/_4332_ ), .CK(clock ), .Q(\RegFile/reg_2 [26] ), .QN(\RegFile/_4151_ ) );
DFF_X1 \RegFile/_7954_ ( .D(\RegFile/_4333_ ), .CK(clock ), .Q(\RegFile/reg_2 [27] ), .QN(\RegFile/_4150_ ) );
DFF_X1 \RegFile/_7955_ ( .D(\RegFile/_4334_ ), .CK(clock ), .Q(\RegFile/reg_2 [28] ), .QN(\RegFile/_4149_ ) );
DFF_X1 \RegFile/_7956_ ( .D(\RegFile/_4335_ ), .CK(clock ), .Q(\RegFile/reg_2 [29] ), .QN(\RegFile/_4148_ ) );
DFF_X1 \RegFile/_7957_ ( .D(\RegFile/_4336_ ), .CK(clock ), .Q(\RegFile/reg_2 [30] ), .QN(\RegFile/_4147_ ) );
DFF_X1 \RegFile/_7958_ ( .D(\RegFile/_4337_ ), .CK(clock ), .Q(\RegFile/reg_2 [31] ), .QN(\RegFile/_4146_ ) );
DFF_X1 \RegFile/_7959_ ( .D(\RegFile/_4338_ ), .CK(clock ), .Q(\RegFile/reg_3 [0] ), .QN(\RegFile/_4145_ ) );
DFF_X1 \RegFile/_7960_ ( .D(\RegFile/_4339_ ), .CK(clock ), .Q(\RegFile/reg_3 [1] ), .QN(\RegFile/_4144_ ) );
DFF_X1 \RegFile/_7961_ ( .D(\RegFile/_4340_ ), .CK(clock ), .Q(\RegFile/reg_3 [2] ), .QN(\RegFile/_4143_ ) );
DFF_X1 \RegFile/_7962_ ( .D(\RegFile/_4341_ ), .CK(clock ), .Q(\RegFile/reg_3 [3] ), .QN(\RegFile/_4142_ ) );
DFF_X1 \RegFile/_7963_ ( .D(\RegFile/_4342_ ), .CK(clock ), .Q(\RegFile/reg_3 [4] ), .QN(\RegFile/_4141_ ) );
DFF_X1 \RegFile/_7964_ ( .D(\RegFile/_4343_ ), .CK(clock ), .Q(\RegFile/reg_3 [5] ), .QN(\RegFile/_4140_ ) );
DFF_X1 \RegFile/_7965_ ( .D(\RegFile/_4344_ ), .CK(clock ), .Q(\RegFile/reg_3 [6] ), .QN(\RegFile/_4139_ ) );
DFF_X1 \RegFile/_7966_ ( .D(\RegFile/_4345_ ), .CK(clock ), .Q(\RegFile/reg_3 [7] ), .QN(\RegFile/_4138_ ) );
DFF_X1 \RegFile/_7967_ ( .D(\RegFile/_4346_ ), .CK(clock ), .Q(\RegFile/reg_3 [8] ), .QN(\RegFile/_4137_ ) );
DFF_X1 \RegFile/_7968_ ( .D(\RegFile/_4347_ ), .CK(clock ), .Q(\RegFile/reg_3 [9] ), .QN(\RegFile/_4136_ ) );
DFF_X1 \RegFile/_7969_ ( .D(\RegFile/_4348_ ), .CK(clock ), .Q(\RegFile/reg_3 [10] ), .QN(\RegFile/_4135_ ) );
DFF_X1 \RegFile/_7970_ ( .D(\RegFile/_4349_ ), .CK(clock ), .Q(\RegFile/reg_3 [11] ), .QN(\RegFile/_4134_ ) );
DFF_X1 \RegFile/_7971_ ( .D(\RegFile/_4350_ ), .CK(clock ), .Q(\RegFile/reg_3 [12] ), .QN(\RegFile/_4133_ ) );
DFF_X1 \RegFile/_7972_ ( .D(\RegFile/_4351_ ), .CK(clock ), .Q(\RegFile/reg_3 [13] ), .QN(\RegFile/_4132_ ) );
DFF_X1 \RegFile/_7973_ ( .D(\RegFile/_4352_ ), .CK(clock ), .Q(\RegFile/reg_3 [14] ), .QN(\RegFile/_4131_ ) );
DFF_X1 \RegFile/_7974_ ( .D(\RegFile/_4353_ ), .CK(clock ), .Q(\RegFile/reg_3 [15] ), .QN(\RegFile/_4130_ ) );
DFF_X1 \RegFile/_7975_ ( .D(\RegFile/_4354_ ), .CK(clock ), .Q(\RegFile/reg_3 [16] ), .QN(\RegFile/_4129_ ) );
DFF_X1 \RegFile/_7976_ ( .D(\RegFile/_4355_ ), .CK(clock ), .Q(\RegFile/reg_3 [17] ), .QN(\RegFile/_4128_ ) );
DFF_X1 \RegFile/_7977_ ( .D(\RegFile/_4356_ ), .CK(clock ), .Q(\RegFile/reg_3 [18] ), .QN(\RegFile/_4127_ ) );
DFF_X1 \RegFile/_7978_ ( .D(\RegFile/_4357_ ), .CK(clock ), .Q(\RegFile/reg_3 [19] ), .QN(\RegFile/_4126_ ) );
DFF_X1 \RegFile/_7979_ ( .D(\RegFile/_4358_ ), .CK(clock ), .Q(\RegFile/reg_3 [20] ), .QN(\RegFile/_4125_ ) );
DFF_X1 \RegFile/_7980_ ( .D(\RegFile/_4359_ ), .CK(clock ), .Q(\RegFile/reg_3 [21] ), .QN(\RegFile/_4124_ ) );
DFF_X1 \RegFile/_7981_ ( .D(\RegFile/_4360_ ), .CK(clock ), .Q(\RegFile/reg_3 [22] ), .QN(\RegFile/_4123_ ) );
DFF_X1 \RegFile/_7982_ ( .D(\RegFile/_4361_ ), .CK(clock ), .Q(\RegFile/reg_3 [23] ), .QN(\RegFile/_4122_ ) );
DFF_X1 \RegFile/_7983_ ( .D(\RegFile/_4362_ ), .CK(clock ), .Q(\RegFile/reg_3 [24] ), .QN(\RegFile/_4121_ ) );
DFF_X1 \RegFile/_7984_ ( .D(\RegFile/_4363_ ), .CK(clock ), .Q(\RegFile/reg_3 [25] ), .QN(\RegFile/_4120_ ) );
DFF_X1 \RegFile/_7985_ ( .D(\RegFile/_4364_ ), .CK(clock ), .Q(\RegFile/reg_3 [26] ), .QN(\RegFile/_4119_ ) );
DFF_X1 \RegFile/_7986_ ( .D(\RegFile/_4365_ ), .CK(clock ), .Q(\RegFile/reg_3 [27] ), .QN(\RegFile/_4118_ ) );
DFF_X1 \RegFile/_7987_ ( .D(\RegFile/_4366_ ), .CK(clock ), .Q(\RegFile/reg_3 [28] ), .QN(\RegFile/_4117_ ) );
DFF_X1 \RegFile/_7988_ ( .D(\RegFile/_4367_ ), .CK(clock ), .Q(\RegFile/reg_3 [29] ), .QN(\RegFile/_4116_ ) );
DFF_X1 \RegFile/_7989_ ( .D(\RegFile/_4368_ ), .CK(clock ), .Q(\RegFile/reg_3 [30] ), .QN(\RegFile/_4115_ ) );
DFF_X1 \RegFile/_7990_ ( .D(\RegFile/_4369_ ), .CK(clock ), .Q(\RegFile/reg_3 [31] ), .QN(\RegFile/_4114_ ) );
DFF_X1 \RegFile/_7991_ ( .D(\RegFile/_4370_ ), .CK(clock ), .Q(\RegFile/reg_4 [0] ), .QN(\RegFile/_4113_ ) );
DFF_X1 \RegFile/_7992_ ( .D(\RegFile/_4371_ ), .CK(clock ), .Q(\RegFile/reg_4 [1] ), .QN(\RegFile/_4112_ ) );
DFF_X1 \RegFile/_7993_ ( .D(\RegFile/_4372_ ), .CK(clock ), .Q(\RegFile/reg_4 [2] ), .QN(\RegFile/_4111_ ) );
DFF_X1 \RegFile/_7994_ ( .D(\RegFile/_4373_ ), .CK(clock ), .Q(\RegFile/reg_4 [3] ), .QN(\RegFile/_4110_ ) );
DFF_X1 \RegFile/_7995_ ( .D(\RegFile/_4374_ ), .CK(clock ), .Q(\RegFile/reg_4 [4] ), .QN(\RegFile/_4109_ ) );
DFF_X1 \RegFile/_7996_ ( .D(\RegFile/_4375_ ), .CK(clock ), .Q(\RegFile/reg_4 [5] ), .QN(\RegFile/_4108_ ) );
DFF_X1 \RegFile/_7997_ ( .D(\RegFile/_4376_ ), .CK(clock ), .Q(\RegFile/reg_4 [6] ), .QN(\RegFile/_4107_ ) );
DFF_X1 \RegFile/_7998_ ( .D(\RegFile/_4377_ ), .CK(clock ), .Q(\RegFile/reg_4 [7] ), .QN(\RegFile/_4106_ ) );
DFF_X1 \RegFile/_7999_ ( .D(\RegFile/_4378_ ), .CK(clock ), .Q(\RegFile/reg_4 [8] ), .QN(\RegFile/_4105_ ) );
DFF_X1 \RegFile/_8000_ ( .D(\RegFile/_4379_ ), .CK(clock ), .Q(\RegFile/reg_4 [9] ), .QN(\RegFile/_4104_ ) );
DFF_X1 \RegFile/_8001_ ( .D(\RegFile/_4380_ ), .CK(clock ), .Q(\RegFile/reg_4 [10] ), .QN(\RegFile/_4103_ ) );
DFF_X1 \RegFile/_8002_ ( .D(\RegFile/_4381_ ), .CK(clock ), .Q(\RegFile/reg_4 [11] ), .QN(\RegFile/_4102_ ) );
DFF_X1 \RegFile/_8003_ ( .D(\RegFile/_4382_ ), .CK(clock ), .Q(\RegFile/reg_4 [12] ), .QN(\RegFile/_4101_ ) );
DFF_X1 \RegFile/_8004_ ( .D(\RegFile/_4383_ ), .CK(clock ), .Q(\RegFile/reg_4 [13] ), .QN(\RegFile/_4100_ ) );
DFF_X1 \RegFile/_8005_ ( .D(\RegFile/_4384_ ), .CK(clock ), .Q(\RegFile/reg_4 [14] ), .QN(\RegFile/_4099_ ) );
DFF_X1 \RegFile/_8006_ ( .D(\RegFile/_4385_ ), .CK(clock ), .Q(\RegFile/reg_4 [15] ), .QN(\RegFile/_4098_ ) );
DFF_X1 \RegFile/_8007_ ( .D(\RegFile/_4386_ ), .CK(clock ), .Q(\RegFile/reg_4 [16] ), .QN(\RegFile/_4097_ ) );
DFF_X1 \RegFile/_8008_ ( .D(\RegFile/_4387_ ), .CK(clock ), .Q(\RegFile/reg_4 [17] ), .QN(\RegFile/_4096_ ) );
DFF_X1 \RegFile/_8009_ ( .D(\RegFile/_4388_ ), .CK(clock ), .Q(\RegFile/reg_4 [18] ), .QN(\RegFile/_4095_ ) );
DFF_X1 \RegFile/_8010_ ( .D(\RegFile/_4389_ ), .CK(clock ), .Q(\RegFile/reg_4 [19] ), .QN(\RegFile/_4094_ ) );
DFF_X1 \RegFile/_8011_ ( .D(\RegFile/_4390_ ), .CK(clock ), .Q(\RegFile/reg_4 [20] ), .QN(\RegFile/_4093_ ) );
DFF_X1 \RegFile/_8012_ ( .D(\RegFile/_4391_ ), .CK(clock ), .Q(\RegFile/reg_4 [21] ), .QN(\RegFile/_4092_ ) );
DFF_X1 \RegFile/_8013_ ( .D(\RegFile/_4392_ ), .CK(clock ), .Q(\RegFile/reg_4 [22] ), .QN(\RegFile/_4091_ ) );
DFF_X1 \RegFile/_8014_ ( .D(\RegFile/_4393_ ), .CK(clock ), .Q(\RegFile/reg_4 [23] ), .QN(\RegFile/_4090_ ) );
DFF_X1 \RegFile/_8015_ ( .D(\RegFile/_4394_ ), .CK(clock ), .Q(\RegFile/reg_4 [24] ), .QN(\RegFile/_4089_ ) );
DFF_X1 \RegFile/_8016_ ( .D(\RegFile/_4395_ ), .CK(clock ), .Q(\RegFile/reg_4 [25] ), .QN(\RegFile/_4088_ ) );
DFF_X1 \RegFile/_8017_ ( .D(\RegFile/_4396_ ), .CK(clock ), .Q(\RegFile/reg_4 [26] ), .QN(\RegFile/_4087_ ) );
DFF_X1 \RegFile/_8018_ ( .D(\RegFile/_4397_ ), .CK(clock ), .Q(\RegFile/reg_4 [27] ), .QN(\RegFile/_4086_ ) );
DFF_X1 \RegFile/_8019_ ( .D(\RegFile/_4398_ ), .CK(clock ), .Q(\RegFile/reg_4 [28] ), .QN(\RegFile/_4085_ ) );
DFF_X1 \RegFile/_8020_ ( .D(\RegFile/_4399_ ), .CK(clock ), .Q(\RegFile/reg_4 [29] ), .QN(\RegFile/_4084_ ) );
DFF_X1 \RegFile/_8021_ ( .D(\RegFile/_4400_ ), .CK(clock ), .Q(\RegFile/reg_4 [30] ), .QN(\RegFile/_4083_ ) );
DFF_X1 \RegFile/_8022_ ( .D(\RegFile/_4401_ ), .CK(clock ), .Q(\RegFile/reg_4 [31] ), .QN(\RegFile/_4082_ ) );
DFF_X1 \RegFile/_8023_ ( .D(\RegFile/_4402_ ), .CK(clock ), .Q(\RegFile/reg_5 [0] ), .QN(\RegFile/_4081_ ) );
DFF_X1 \RegFile/_8024_ ( .D(\RegFile/_4403_ ), .CK(clock ), .Q(\RegFile/reg_5 [1] ), .QN(\RegFile/_4080_ ) );
DFF_X1 \RegFile/_8025_ ( .D(\RegFile/_4404_ ), .CK(clock ), .Q(\RegFile/reg_5 [2] ), .QN(\RegFile/_4079_ ) );
DFF_X1 \RegFile/_8026_ ( .D(\RegFile/_4405_ ), .CK(clock ), .Q(\RegFile/reg_5 [3] ), .QN(\RegFile/_4078_ ) );
DFF_X1 \RegFile/_8027_ ( .D(\RegFile/_4406_ ), .CK(clock ), .Q(\RegFile/reg_5 [4] ), .QN(\RegFile/_4077_ ) );
DFF_X1 \RegFile/_8028_ ( .D(\RegFile/_4407_ ), .CK(clock ), .Q(\RegFile/reg_5 [5] ), .QN(\RegFile/_4076_ ) );
DFF_X1 \RegFile/_8029_ ( .D(\RegFile/_4408_ ), .CK(clock ), .Q(\RegFile/reg_5 [6] ), .QN(\RegFile/_4075_ ) );
DFF_X1 \RegFile/_8030_ ( .D(\RegFile/_4409_ ), .CK(clock ), .Q(\RegFile/reg_5 [7] ), .QN(\RegFile/_4074_ ) );
DFF_X1 \RegFile/_8031_ ( .D(\RegFile/_4410_ ), .CK(clock ), .Q(\RegFile/reg_5 [8] ), .QN(\RegFile/_4073_ ) );
DFF_X1 \RegFile/_8032_ ( .D(\RegFile/_4411_ ), .CK(clock ), .Q(\RegFile/reg_5 [9] ), .QN(\RegFile/_4072_ ) );
DFF_X1 \RegFile/_8033_ ( .D(\RegFile/_4412_ ), .CK(clock ), .Q(\RegFile/reg_5 [10] ), .QN(\RegFile/_4071_ ) );
DFF_X1 \RegFile/_8034_ ( .D(\RegFile/_4413_ ), .CK(clock ), .Q(\RegFile/reg_5 [11] ), .QN(\RegFile/_4070_ ) );
DFF_X1 \RegFile/_8035_ ( .D(\RegFile/_4414_ ), .CK(clock ), .Q(\RegFile/reg_5 [12] ), .QN(\RegFile/_4069_ ) );
DFF_X1 \RegFile/_8036_ ( .D(\RegFile/_4415_ ), .CK(clock ), .Q(\RegFile/reg_5 [13] ), .QN(\RegFile/_4068_ ) );
DFF_X1 \RegFile/_8037_ ( .D(\RegFile/_4416_ ), .CK(clock ), .Q(\RegFile/reg_5 [14] ), .QN(\RegFile/_4067_ ) );
DFF_X1 \RegFile/_8038_ ( .D(\RegFile/_4417_ ), .CK(clock ), .Q(\RegFile/reg_5 [15] ), .QN(\RegFile/_4066_ ) );
DFF_X1 \RegFile/_8039_ ( .D(\RegFile/_4418_ ), .CK(clock ), .Q(\RegFile/reg_5 [16] ), .QN(\RegFile/_4065_ ) );
DFF_X1 \RegFile/_8040_ ( .D(\RegFile/_4419_ ), .CK(clock ), .Q(\RegFile/reg_5 [17] ), .QN(\RegFile/_4064_ ) );
DFF_X1 \RegFile/_8041_ ( .D(\RegFile/_4420_ ), .CK(clock ), .Q(\RegFile/reg_5 [18] ), .QN(\RegFile/_4063_ ) );
DFF_X1 \RegFile/_8042_ ( .D(\RegFile/_4421_ ), .CK(clock ), .Q(\RegFile/reg_5 [19] ), .QN(\RegFile/_4062_ ) );
DFF_X1 \RegFile/_8043_ ( .D(\RegFile/_4422_ ), .CK(clock ), .Q(\RegFile/reg_5 [20] ), .QN(\RegFile/_4061_ ) );
DFF_X1 \RegFile/_8044_ ( .D(\RegFile/_4423_ ), .CK(clock ), .Q(\RegFile/reg_5 [21] ), .QN(\RegFile/_4060_ ) );
DFF_X1 \RegFile/_8045_ ( .D(\RegFile/_4424_ ), .CK(clock ), .Q(\RegFile/reg_5 [22] ), .QN(\RegFile/_4059_ ) );
DFF_X1 \RegFile/_8046_ ( .D(\RegFile/_4425_ ), .CK(clock ), .Q(\RegFile/reg_5 [23] ), .QN(\RegFile/_4058_ ) );
DFF_X1 \RegFile/_8047_ ( .D(\RegFile/_4426_ ), .CK(clock ), .Q(\RegFile/reg_5 [24] ), .QN(\RegFile/_4057_ ) );
DFF_X1 \RegFile/_8048_ ( .D(\RegFile/_4427_ ), .CK(clock ), .Q(\RegFile/reg_5 [25] ), .QN(\RegFile/_4056_ ) );
DFF_X1 \RegFile/_8049_ ( .D(\RegFile/_4428_ ), .CK(clock ), .Q(\RegFile/reg_5 [26] ), .QN(\RegFile/_4055_ ) );
DFF_X1 \RegFile/_8050_ ( .D(\RegFile/_4429_ ), .CK(clock ), .Q(\RegFile/reg_5 [27] ), .QN(\RegFile/_4054_ ) );
DFF_X1 \RegFile/_8051_ ( .D(\RegFile/_4430_ ), .CK(clock ), .Q(\RegFile/reg_5 [28] ), .QN(\RegFile/_4053_ ) );
DFF_X1 \RegFile/_8052_ ( .D(\RegFile/_4431_ ), .CK(clock ), .Q(\RegFile/reg_5 [29] ), .QN(\RegFile/_4052_ ) );
DFF_X1 \RegFile/_8053_ ( .D(\RegFile/_4432_ ), .CK(clock ), .Q(\RegFile/reg_5 [30] ), .QN(\RegFile/_4051_ ) );
DFF_X1 \RegFile/_8054_ ( .D(\RegFile/_4433_ ), .CK(clock ), .Q(\RegFile/reg_5 [31] ), .QN(\RegFile/_4050_ ) );
DFF_X1 \RegFile/_8055_ ( .D(\RegFile/_4434_ ), .CK(clock ), .Q(\RegFile/reg_6 [0] ), .QN(\RegFile/_4049_ ) );
DFF_X1 \RegFile/_8056_ ( .D(\RegFile/_4435_ ), .CK(clock ), .Q(\RegFile/reg_6 [1] ), .QN(\RegFile/_4048_ ) );
DFF_X1 \RegFile/_8057_ ( .D(\RegFile/_4436_ ), .CK(clock ), .Q(\RegFile/reg_6 [2] ), .QN(\RegFile/_4047_ ) );
DFF_X1 \RegFile/_8058_ ( .D(\RegFile/_4437_ ), .CK(clock ), .Q(\RegFile/reg_6 [3] ), .QN(\RegFile/_4046_ ) );
DFF_X1 \RegFile/_8059_ ( .D(\RegFile/_4438_ ), .CK(clock ), .Q(\RegFile/reg_6 [4] ), .QN(\RegFile/_4045_ ) );
DFF_X1 \RegFile/_8060_ ( .D(\RegFile/_4439_ ), .CK(clock ), .Q(\RegFile/reg_6 [5] ), .QN(\RegFile/_4044_ ) );
DFF_X1 \RegFile/_8061_ ( .D(\RegFile/_4440_ ), .CK(clock ), .Q(\RegFile/reg_6 [6] ), .QN(\RegFile/_4043_ ) );
DFF_X1 \RegFile/_8062_ ( .D(\RegFile/_4441_ ), .CK(clock ), .Q(\RegFile/reg_6 [7] ), .QN(\RegFile/_4042_ ) );
DFF_X1 \RegFile/_8063_ ( .D(\RegFile/_4442_ ), .CK(clock ), .Q(\RegFile/reg_6 [8] ), .QN(\RegFile/_4041_ ) );
DFF_X1 \RegFile/_8064_ ( .D(\RegFile/_4443_ ), .CK(clock ), .Q(\RegFile/reg_6 [9] ), .QN(\RegFile/_4040_ ) );
DFF_X1 \RegFile/_8065_ ( .D(\RegFile/_4444_ ), .CK(clock ), .Q(\RegFile/reg_6 [10] ), .QN(\RegFile/_4039_ ) );
DFF_X1 \RegFile/_8066_ ( .D(\RegFile/_4445_ ), .CK(clock ), .Q(\RegFile/reg_6 [11] ), .QN(\RegFile/_4038_ ) );
DFF_X1 \RegFile/_8067_ ( .D(\RegFile/_4446_ ), .CK(clock ), .Q(\RegFile/reg_6 [12] ), .QN(\RegFile/_4037_ ) );
DFF_X1 \RegFile/_8068_ ( .D(\RegFile/_4447_ ), .CK(clock ), .Q(\RegFile/reg_6 [13] ), .QN(\RegFile/_4036_ ) );
DFF_X1 \RegFile/_8069_ ( .D(\RegFile/_4448_ ), .CK(clock ), .Q(\RegFile/reg_6 [14] ), .QN(\RegFile/_4035_ ) );
DFF_X1 \RegFile/_8070_ ( .D(\RegFile/_4449_ ), .CK(clock ), .Q(\RegFile/reg_6 [15] ), .QN(\RegFile/_4034_ ) );
DFF_X1 \RegFile/_8071_ ( .D(\RegFile/_4450_ ), .CK(clock ), .Q(\RegFile/reg_6 [16] ), .QN(\RegFile/_4033_ ) );
DFF_X1 \RegFile/_8072_ ( .D(\RegFile/_4451_ ), .CK(clock ), .Q(\RegFile/reg_6 [17] ), .QN(\RegFile/_4032_ ) );
DFF_X1 \RegFile/_8073_ ( .D(\RegFile/_4452_ ), .CK(clock ), .Q(\RegFile/reg_6 [18] ), .QN(\RegFile/_4031_ ) );
DFF_X1 \RegFile/_8074_ ( .D(\RegFile/_4453_ ), .CK(clock ), .Q(\RegFile/reg_6 [19] ), .QN(\RegFile/_4030_ ) );
DFF_X1 \RegFile/_8075_ ( .D(\RegFile/_4454_ ), .CK(clock ), .Q(\RegFile/reg_6 [20] ), .QN(\RegFile/_4029_ ) );
DFF_X1 \RegFile/_8076_ ( .D(\RegFile/_4455_ ), .CK(clock ), .Q(\RegFile/reg_6 [21] ), .QN(\RegFile/_4028_ ) );
DFF_X1 \RegFile/_8077_ ( .D(\RegFile/_4456_ ), .CK(clock ), .Q(\RegFile/reg_6 [22] ), .QN(\RegFile/_4027_ ) );
DFF_X1 \RegFile/_8078_ ( .D(\RegFile/_4457_ ), .CK(clock ), .Q(\RegFile/reg_6 [23] ), .QN(\RegFile/_4026_ ) );
DFF_X1 \RegFile/_8079_ ( .D(\RegFile/_4458_ ), .CK(clock ), .Q(\RegFile/reg_6 [24] ), .QN(\RegFile/_4025_ ) );
DFF_X1 \RegFile/_8080_ ( .D(\RegFile/_4459_ ), .CK(clock ), .Q(\RegFile/reg_6 [25] ), .QN(\RegFile/_4024_ ) );
DFF_X1 \RegFile/_8081_ ( .D(\RegFile/_4460_ ), .CK(clock ), .Q(\RegFile/reg_6 [26] ), .QN(\RegFile/_4023_ ) );
DFF_X1 \RegFile/_8082_ ( .D(\RegFile/_4461_ ), .CK(clock ), .Q(\RegFile/reg_6 [27] ), .QN(\RegFile/_4022_ ) );
DFF_X1 \RegFile/_8083_ ( .D(\RegFile/_4462_ ), .CK(clock ), .Q(\RegFile/reg_6 [28] ), .QN(\RegFile/_4021_ ) );
DFF_X1 \RegFile/_8084_ ( .D(\RegFile/_4463_ ), .CK(clock ), .Q(\RegFile/reg_6 [29] ), .QN(\RegFile/_4020_ ) );
DFF_X1 \RegFile/_8085_ ( .D(\RegFile/_4464_ ), .CK(clock ), .Q(\RegFile/reg_6 [30] ), .QN(\RegFile/_4019_ ) );
DFF_X1 \RegFile/_8086_ ( .D(\RegFile/_4465_ ), .CK(clock ), .Q(\RegFile/reg_6 [31] ), .QN(\RegFile/_4018_ ) );
DFF_X1 \RegFile/_8087_ ( .D(\RegFile/_4466_ ), .CK(clock ), .Q(\RegFile/reg_7 [0] ), .QN(\RegFile/_4017_ ) );
DFF_X1 \RegFile/_8088_ ( .D(\RegFile/_4467_ ), .CK(clock ), .Q(\RegFile/reg_7 [1] ), .QN(\RegFile/_4016_ ) );
DFF_X1 \RegFile/_8089_ ( .D(\RegFile/_4468_ ), .CK(clock ), .Q(\RegFile/reg_7 [2] ), .QN(\RegFile/_4015_ ) );
DFF_X1 \RegFile/_8090_ ( .D(\RegFile/_4469_ ), .CK(clock ), .Q(\RegFile/reg_7 [3] ), .QN(\RegFile/_4014_ ) );
DFF_X1 \RegFile/_8091_ ( .D(\RegFile/_4470_ ), .CK(clock ), .Q(\RegFile/reg_7 [4] ), .QN(\RegFile/_4013_ ) );
DFF_X1 \RegFile/_8092_ ( .D(\RegFile/_4471_ ), .CK(clock ), .Q(\RegFile/reg_7 [5] ), .QN(\RegFile/_4012_ ) );
DFF_X1 \RegFile/_8093_ ( .D(\RegFile/_4472_ ), .CK(clock ), .Q(\RegFile/reg_7 [6] ), .QN(\RegFile/_4011_ ) );
DFF_X1 \RegFile/_8094_ ( .D(\RegFile/_4473_ ), .CK(clock ), .Q(\RegFile/reg_7 [7] ), .QN(\RegFile/_4010_ ) );
DFF_X1 \RegFile/_8095_ ( .D(\RegFile/_4474_ ), .CK(clock ), .Q(\RegFile/reg_7 [8] ), .QN(\RegFile/_4009_ ) );
DFF_X1 \RegFile/_8096_ ( .D(\RegFile/_4475_ ), .CK(clock ), .Q(\RegFile/reg_7 [9] ), .QN(\RegFile/_4008_ ) );
DFF_X1 \RegFile/_8097_ ( .D(\RegFile/_4476_ ), .CK(clock ), .Q(\RegFile/reg_7 [10] ), .QN(\RegFile/_4007_ ) );
DFF_X1 \RegFile/_8098_ ( .D(\RegFile/_4477_ ), .CK(clock ), .Q(\RegFile/reg_7 [11] ), .QN(\RegFile/_4006_ ) );
DFF_X1 \RegFile/_8099_ ( .D(\RegFile/_4478_ ), .CK(clock ), .Q(\RegFile/reg_7 [12] ), .QN(\RegFile/_4005_ ) );
DFF_X1 \RegFile/_8100_ ( .D(\RegFile/_4479_ ), .CK(clock ), .Q(\RegFile/reg_7 [13] ), .QN(\RegFile/_4004_ ) );
DFF_X1 \RegFile/_8101_ ( .D(\RegFile/_4480_ ), .CK(clock ), .Q(\RegFile/reg_7 [14] ), .QN(\RegFile/_4003_ ) );
DFF_X1 \RegFile/_8102_ ( .D(\RegFile/_4481_ ), .CK(clock ), .Q(\RegFile/reg_7 [15] ), .QN(\RegFile/_4002_ ) );
DFF_X1 \RegFile/_8103_ ( .D(\RegFile/_4482_ ), .CK(clock ), .Q(\RegFile/reg_7 [16] ), .QN(\RegFile/_4001_ ) );
DFF_X1 \RegFile/_8104_ ( .D(\RegFile/_4483_ ), .CK(clock ), .Q(\RegFile/reg_7 [17] ), .QN(\RegFile/_4000_ ) );
DFF_X1 \RegFile/_8105_ ( .D(\RegFile/_4484_ ), .CK(clock ), .Q(\RegFile/reg_7 [18] ), .QN(\RegFile/_3999_ ) );
DFF_X1 \RegFile/_8106_ ( .D(\RegFile/_4485_ ), .CK(clock ), .Q(\RegFile/reg_7 [19] ), .QN(\RegFile/_3998_ ) );
DFF_X1 \RegFile/_8107_ ( .D(\RegFile/_4486_ ), .CK(clock ), .Q(\RegFile/reg_7 [20] ), .QN(\RegFile/_3997_ ) );
DFF_X1 \RegFile/_8108_ ( .D(\RegFile/_4487_ ), .CK(clock ), .Q(\RegFile/reg_7 [21] ), .QN(\RegFile/_3996_ ) );
DFF_X1 \RegFile/_8109_ ( .D(\RegFile/_4488_ ), .CK(clock ), .Q(\RegFile/reg_7 [22] ), .QN(\RegFile/_3995_ ) );
DFF_X1 \RegFile/_8110_ ( .D(\RegFile/_4489_ ), .CK(clock ), .Q(\RegFile/reg_7 [23] ), .QN(\RegFile/_3994_ ) );
DFF_X1 \RegFile/_8111_ ( .D(\RegFile/_4490_ ), .CK(clock ), .Q(\RegFile/reg_7 [24] ), .QN(\RegFile/_3993_ ) );
DFF_X1 \RegFile/_8112_ ( .D(\RegFile/_4491_ ), .CK(clock ), .Q(\RegFile/reg_7 [25] ), .QN(\RegFile/_3992_ ) );
DFF_X1 \RegFile/_8113_ ( .D(\RegFile/_4492_ ), .CK(clock ), .Q(\RegFile/reg_7 [26] ), .QN(\RegFile/_3991_ ) );
DFF_X1 \RegFile/_8114_ ( .D(\RegFile/_4493_ ), .CK(clock ), .Q(\RegFile/reg_7 [27] ), .QN(\RegFile/_3990_ ) );
DFF_X1 \RegFile/_8115_ ( .D(\RegFile/_4494_ ), .CK(clock ), .Q(\RegFile/reg_7 [28] ), .QN(\RegFile/_3989_ ) );
DFF_X1 \RegFile/_8116_ ( .D(\RegFile/_4495_ ), .CK(clock ), .Q(\RegFile/reg_7 [29] ), .QN(\RegFile/_3988_ ) );
DFF_X1 \RegFile/_8117_ ( .D(\RegFile/_4496_ ), .CK(clock ), .Q(\RegFile/reg_7 [30] ), .QN(\RegFile/_3987_ ) );
DFF_X1 \RegFile/_8118_ ( .D(\RegFile/_4497_ ), .CK(clock ), .Q(\RegFile/reg_7 [31] ), .QN(\RegFile/_3986_ ) );
DFF_X1 \RegFile/_8119_ ( .D(\RegFile/_4498_ ), .CK(clock ), .Q(\RegFile/reg_8 [0] ), .QN(\RegFile/_3985_ ) );
DFF_X1 \RegFile/_8120_ ( .D(\RegFile/_4499_ ), .CK(clock ), .Q(\RegFile/reg_8 [1] ), .QN(\RegFile/_3984_ ) );
DFF_X1 \RegFile/_8121_ ( .D(\RegFile/_4500_ ), .CK(clock ), .Q(\RegFile/reg_8 [2] ), .QN(\RegFile/_3983_ ) );
DFF_X1 \RegFile/_8122_ ( .D(\RegFile/_4501_ ), .CK(clock ), .Q(\RegFile/reg_8 [3] ), .QN(\RegFile/_3982_ ) );
DFF_X1 \RegFile/_8123_ ( .D(\RegFile/_4502_ ), .CK(clock ), .Q(\RegFile/reg_8 [4] ), .QN(\RegFile/_3981_ ) );
DFF_X1 \RegFile/_8124_ ( .D(\RegFile/_4503_ ), .CK(clock ), .Q(\RegFile/reg_8 [5] ), .QN(\RegFile/_3980_ ) );
DFF_X1 \RegFile/_8125_ ( .D(\RegFile/_4504_ ), .CK(clock ), .Q(\RegFile/reg_8 [6] ), .QN(\RegFile/_3979_ ) );
DFF_X1 \RegFile/_8126_ ( .D(\RegFile/_4505_ ), .CK(clock ), .Q(\RegFile/reg_8 [7] ), .QN(\RegFile/_3978_ ) );
DFF_X1 \RegFile/_8127_ ( .D(\RegFile/_4506_ ), .CK(clock ), .Q(\RegFile/reg_8 [8] ), .QN(\RegFile/_3977_ ) );
DFF_X1 \RegFile/_8128_ ( .D(\RegFile/_4507_ ), .CK(clock ), .Q(\RegFile/reg_8 [9] ), .QN(\RegFile/_3976_ ) );
DFF_X1 \RegFile/_8129_ ( .D(\RegFile/_4508_ ), .CK(clock ), .Q(\RegFile/reg_8 [10] ), .QN(\RegFile/_3975_ ) );
DFF_X1 \RegFile/_8130_ ( .D(\RegFile/_4509_ ), .CK(clock ), .Q(\RegFile/reg_8 [11] ), .QN(\RegFile/_3974_ ) );
DFF_X1 \RegFile/_8131_ ( .D(\RegFile/_4510_ ), .CK(clock ), .Q(\RegFile/reg_8 [12] ), .QN(\RegFile/_3973_ ) );
DFF_X1 \RegFile/_8132_ ( .D(\RegFile/_4511_ ), .CK(clock ), .Q(\RegFile/reg_8 [13] ), .QN(\RegFile/_3972_ ) );
DFF_X1 \RegFile/_8133_ ( .D(\RegFile/_4512_ ), .CK(clock ), .Q(\RegFile/reg_8 [14] ), .QN(\RegFile/_3971_ ) );
DFF_X1 \RegFile/_8134_ ( .D(\RegFile/_4513_ ), .CK(clock ), .Q(\RegFile/reg_8 [15] ), .QN(\RegFile/_3970_ ) );
DFF_X1 \RegFile/_8135_ ( .D(\RegFile/_4514_ ), .CK(clock ), .Q(\RegFile/reg_8 [16] ), .QN(\RegFile/_3969_ ) );
DFF_X1 \RegFile/_8136_ ( .D(\RegFile/_4515_ ), .CK(clock ), .Q(\RegFile/reg_8 [17] ), .QN(\RegFile/_3968_ ) );
DFF_X1 \RegFile/_8137_ ( .D(\RegFile/_4516_ ), .CK(clock ), .Q(\RegFile/reg_8 [18] ), .QN(\RegFile/_3967_ ) );
DFF_X1 \RegFile/_8138_ ( .D(\RegFile/_4517_ ), .CK(clock ), .Q(\RegFile/reg_8 [19] ), .QN(\RegFile/_3966_ ) );
DFF_X1 \RegFile/_8139_ ( .D(\RegFile/_4518_ ), .CK(clock ), .Q(\RegFile/reg_8 [20] ), .QN(\RegFile/_3965_ ) );
DFF_X1 \RegFile/_8140_ ( .D(\RegFile/_4519_ ), .CK(clock ), .Q(\RegFile/reg_8 [21] ), .QN(\RegFile/_3964_ ) );
DFF_X1 \RegFile/_8141_ ( .D(\RegFile/_4520_ ), .CK(clock ), .Q(\RegFile/reg_8 [22] ), .QN(\RegFile/_3963_ ) );
DFF_X1 \RegFile/_8142_ ( .D(\RegFile/_4521_ ), .CK(clock ), .Q(\RegFile/reg_8 [23] ), .QN(\RegFile/_3962_ ) );
DFF_X1 \RegFile/_8143_ ( .D(\RegFile/_4522_ ), .CK(clock ), .Q(\RegFile/reg_8 [24] ), .QN(\RegFile/_3961_ ) );
DFF_X1 \RegFile/_8144_ ( .D(\RegFile/_4523_ ), .CK(clock ), .Q(\RegFile/reg_8 [25] ), .QN(\RegFile/_3960_ ) );
DFF_X1 \RegFile/_8145_ ( .D(\RegFile/_4524_ ), .CK(clock ), .Q(\RegFile/reg_8 [26] ), .QN(\RegFile/_3959_ ) );
DFF_X1 \RegFile/_8146_ ( .D(\RegFile/_4525_ ), .CK(clock ), .Q(\RegFile/reg_8 [27] ), .QN(\RegFile/_3958_ ) );
DFF_X1 \RegFile/_8147_ ( .D(\RegFile/_4526_ ), .CK(clock ), .Q(\RegFile/reg_8 [28] ), .QN(\RegFile/_3957_ ) );
DFF_X1 \RegFile/_8148_ ( .D(\RegFile/_4527_ ), .CK(clock ), .Q(\RegFile/reg_8 [29] ), .QN(\RegFile/_3956_ ) );
DFF_X1 \RegFile/_8149_ ( .D(\RegFile/_4528_ ), .CK(clock ), .Q(\RegFile/reg_8 [30] ), .QN(\RegFile/_3955_ ) );
DFF_X1 \RegFile/_8150_ ( .D(\RegFile/_4529_ ), .CK(clock ), .Q(\RegFile/reg_8 [31] ), .QN(\RegFile/_3954_ ) );
DFF_X1 \RegFile/_8151_ ( .D(\RegFile/_4530_ ), .CK(clock ), .Q(\RegFile/reg_9 [0] ), .QN(\RegFile/_3953_ ) );
DFF_X1 \RegFile/_8152_ ( .D(\RegFile/_4531_ ), .CK(clock ), .Q(\RegFile/reg_9 [1] ), .QN(\RegFile/_3952_ ) );
DFF_X1 \RegFile/_8153_ ( .D(\RegFile/_4532_ ), .CK(clock ), .Q(\RegFile/reg_9 [2] ), .QN(\RegFile/_3951_ ) );
DFF_X1 \RegFile/_8154_ ( .D(\RegFile/_4533_ ), .CK(clock ), .Q(\RegFile/reg_9 [3] ), .QN(\RegFile/_3950_ ) );
DFF_X1 \RegFile/_8155_ ( .D(\RegFile/_4534_ ), .CK(clock ), .Q(\RegFile/reg_9 [4] ), .QN(\RegFile/_3949_ ) );
DFF_X1 \RegFile/_8156_ ( .D(\RegFile/_4535_ ), .CK(clock ), .Q(\RegFile/reg_9 [5] ), .QN(\RegFile/_3948_ ) );
DFF_X1 \RegFile/_8157_ ( .D(\RegFile/_4536_ ), .CK(clock ), .Q(\RegFile/reg_9 [6] ), .QN(\RegFile/_3947_ ) );
DFF_X1 \RegFile/_8158_ ( .D(\RegFile/_4537_ ), .CK(clock ), .Q(\RegFile/reg_9 [7] ), .QN(\RegFile/_3946_ ) );
DFF_X1 \RegFile/_8159_ ( .D(\RegFile/_4538_ ), .CK(clock ), .Q(\RegFile/reg_9 [8] ), .QN(\RegFile/_3945_ ) );
DFF_X1 \RegFile/_8160_ ( .D(\RegFile/_4539_ ), .CK(clock ), .Q(\RegFile/reg_9 [9] ), .QN(\RegFile/_3944_ ) );
DFF_X1 \RegFile/_8161_ ( .D(\RegFile/_4540_ ), .CK(clock ), .Q(\RegFile/reg_9 [10] ), .QN(\RegFile/_3943_ ) );
DFF_X1 \RegFile/_8162_ ( .D(\RegFile/_4541_ ), .CK(clock ), .Q(\RegFile/reg_9 [11] ), .QN(\RegFile/_3942_ ) );
DFF_X1 \RegFile/_8163_ ( .D(\RegFile/_4542_ ), .CK(clock ), .Q(\RegFile/reg_9 [12] ), .QN(\RegFile/_3941_ ) );
DFF_X1 \RegFile/_8164_ ( .D(\RegFile/_4543_ ), .CK(clock ), .Q(\RegFile/reg_9 [13] ), .QN(\RegFile/_3940_ ) );
DFF_X1 \RegFile/_8165_ ( .D(\RegFile/_4544_ ), .CK(clock ), .Q(\RegFile/reg_9 [14] ), .QN(\RegFile/_3939_ ) );
DFF_X1 \RegFile/_8166_ ( .D(\RegFile/_4545_ ), .CK(clock ), .Q(\RegFile/reg_9 [15] ), .QN(\RegFile/_3938_ ) );
DFF_X1 \RegFile/_8167_ ( .D(\RegFile/_4546_ ), .CK(clock ), .Q(\RegFile/reg_9 [16] ), .QN(\RegFile/_3937_ ) );
DFF_X1 \RegFile/_8168_ ( .D(\RegFile/_4547_ ), .CK(clock ), .Q(\RegFile/reg_9 [17] ), .QN(\RegFile/_3936_ ) );
DFF_X1 \RegFile/_8169_ ( .D(\RegFile/_4548_ ), .CK(clock ), .Q(\RegFile/reg_9 [18] ), .QN(\RegFile/_3935_ ) );
DFF_X1 \RegFile/_8170_ ( .D(\RegFile/_4549_ ), .CK(clock ), .Q(\RegFile/reg_9 [19] ), .QN(\RegFile/_3934_ ) );
DFF_X1 \RegFile/_8171_ ( .D(\RegFile/_4550_ ), .CK(clock ), .Q(\RegFile/reg_9 [20] ), .QN(\RegFile/_3933_ ) );
DFF_X1 \RegFile/_8172_ ( .D(\RegFile/_4551_ ), .CK(clock ), .Q(\RegFile/reg_9 [21] ), .QN(\RegFile/_3932_ ) );
DFF_X1 \RegFile/_8173_ ( .D(\RegFile/_4552_ ), .CK(clock ), .Q(\RegFile/reg_9 [22] ), .QN(\RegFile/_3931_ ) );
DFF_X1 \RegFile/_8174_ ( .D(\RegFile/_4553_ ), .CK(clock ), .Q(\RegFile/reg_9 [23] ), .QN(\RegFile/_3930_ ) );
DFF_X1 \RegFile/_8175_ ( .D(\RegFile/_4554_ ), .CK(clock ), .Q(\RegFile/reg_9 [24] ), .QN(\RegFile/_3929_ ) );
DFF_X1 \RegFile/_8176_ ( .D(\RegFile/_4555_ ), .CK(clock ), .Q(\RegFile/reg_9 [25] ), .QN(\RegFile/_3928_ ) );
DFF_X1 \RegFile/_8177_ ( .D(\RegFile/_4556_ ), .CK(clock ), .Q(\RegFile/reg_9 [26] ), .QN(\RegFile/_3927_ ) );
DFF_X1 \RegFile/_8178_ ( .D(\RegFile/_4557_ ), .CK(clock ), .Q(\RegFile/reg_9 [27] ), .QN(\RegFile/_3926_ ) );
DFF_X1 \RegFile/_8179_ ( .D(\RegFile/_4558_ ), .CK(clock ), .Q(\RegFile/reg_9 [28] ), .QN(\RegFile/_3925_ ) );
DFF_X1 \RegFile/_8180_ ( .D(\RegFile/_4559_ ), .CK(clock ), .Q(\RegFile/reg_9 [29] ), .QN(\RegFile/_3924_ ) );
DFF_X1 \RegFile/_8181_ ( .D(\RegFile/_4560_ ), .CK(clock ), .Q(\RegFile/reg_9 [30] ), .QN(\RegFile/_3923_ ) );
DFF_X1 \RegFile/_8182_ ( .D(\RegFile/_4561_ ), .CK(clock ), .Q(\RegFile/reg_9 [31] ), .QN(\RegFile/_3922_ ) );
DFF_X1 \RegFile/_8183_ ( .D(\RegFile/_4562_ ), .CK(clock ), .Q(\RegFile/reg_10 [0] ), .QN(\RegFile/_3921_ ) );
DFF_X1 \RegFile/_8184_ ( .D(\RegFile/_4563_ ), .CK(clock ), .Q(\RegFile/reg_10 [1] ), .QN(\RegFile/_3920_ ) );
DFF_X1 \RegFile/_8185_ ( .D(\RegFile/_4564_ ), .CK(clock ), .Q(\RegFile/reg_10 [2] ), .QN(\RegFile/_3919_ ) );
DFF_X1 \RegFile/_8186_ ( .D(\RegFile/_4565_ ), .CK(clock ), .Q(\RegFile/reg_10 [3] ), .QN(\RegFile/_3918_ ) );
DFF_X1 \RegFile/_8187_ ( .D(\RegFile/_4566_ ), .CK(clock ), .Q(\RegFile/reg_10 [4] ), .QN(\RegFile/_3917_ ) );
DFF_X1 \RegFile/_8188_ ( .D(\RegFile/_4567_ ), .CK(clock ), .Q(\RegFile/reg_10 [5] ), .QN(\RegFile/_3916_ ) );
DFF_X1 \RegFile/_8189_ ( .D(\RegFile/_4568_ ), .CK(clock ), .Q(\RegFile/reg_10 [6] ), .QN(\RegFile/_3915_ ) );
DFF_X1 \RegFile/_8190_ ( .D(\RegFile/_4569_ ), .CK(clock ), .Q(\RegFile/reg_10 [7] ), .QN(\RegFile/_3914_ ) );
DFF_X1 \RegFile/_8191_ ( .D(\RegFile/_4570_ ), .CK(clock ), .Q(\RegFile/reg_10 [8] ), .QN(\RegFile/_3913_ ) );
DFF_X1 \RegFile/_8192_ ( .D(\RegFile/_4571_ ), .CK(clock ), .Q(\RegFile/reg_10 [9] ), .QN(\RegFile/_3912_ ) );
DFF_X1 \RegFile/_8193_ ( .D(\RegFile/_4572_ ), .CK(clock ), .Q(\RegFile/reg_10 [10] ), .QN(\RegFile/_3911_ ) );
DFF_X1 \RegFile/_8194_ ( .D(\RegFile/_4573_ ), .CK(clock ), .Q(\RegFile/reg_10 [11] ), .QN(\RegFile/_3910_ ) );
DFF_X1 \RegFile/_8195_ ( .D(\RegFile/_4574_ ), .CK(clock ), .Q(\RegFile/reg_10 [12] ), .QN(\RegFile/_3909_ ) );
DFF_X1 \RegFile/_8196_ ( .D(\RegFile/_4575_ ), .CK(clock ), .Q(\RegFile/reg_10 [13] ), .QN(\RegFile/_3908_ ) );
DFF_X1 \RegFile/_8197_ ( .D(\RegFile/_4576_ ), .CK(clock ), .Q(\RegFile/reg_10 [14] ), .QN(\RegFile/_3907_ ) );
DFF_X1 \RegFile/_8198_ ( .D(\RegFile/_4577_ ), .CK(clock ), .Q(\RegFile/reg_10 [15] ), .QN(\RegFile/_3906_ ) );
DFF_X1 \RegFile/_8199_ ( .D(\RegFile/_4578_ ), .CK(clock ), .Q(\RegFile/reg_10 [16] ), .QN(\RegFile/_3905_ ) );
DFF_X1 \RegFile/_8200_ ( .D(\RegFile/_4579_ ), .CK(clock ), .Q(\RegFile/reg_10 [17] ), .QN(\RegFile/_3904_ ) );
DFF_X1 \RegFile/_8201_ ( .D(\RegFile/_4580_ ), .CK(clock ), .Q(\RegFile/reg_10 [18] ), .QN(\RegFile/_3903_ ) );
DFF_X1 \RegFile/_8202_ ( .D(\RegFile/_4581_ ), .CK(clock ), .Q(\RegFile/reg_10 [19] ), .QN(\RegFile/_3902_ ) );
DFF_X1 \RegFile/_8203_ ( .D(\RegFile/_4582_ ), .CK(clock ), .Q(\RegFile/reg_10 [20] ), .QN(\RegFile/_3901_ ) );
DFF_X1 \RegFile/_8204_ ( .D(\RegFile/_4583_ ), .CK(clock ), .Q(\RegFile/reg_10 [21] ), .QN(\RegFile/_3900_ ) );
DFF_X1 \RegFile/_8205_ ( .D(\RegFile/_4584_ ), .CK(clock ), .Q(\RegFile/reg_10 [22] ), .QN(\RegFile/_3899_ ) );
DFF_X1 \RegFile/_8206_ ( .D(\RegFile/_4585_ ), .CK(clock ), .Q(\RegFile/reg_10 [23] ), .QN(\RegFile/_3898_ ) );
DFF_X1 \RegFile/_8207_ ( .D(\RegFile/_4586_ ), .CK(clock ), .Q(\RegFile/reg_10 [24] ), .QN(\RegFile/_3897_ ) );
DFF_X1 \RegFile/_8208_ ( .D(\RegFile/_4587_ ), .CK(clock ), .Q(\RegFile/reg_10 [25] ), .QN(\RegFile/_3896_ ) );
DFF_X1 \RegFile/_8209_ ( .D(\RegFile/_4588_ ), .CK(clock ), .Q(\RegFile/reg_10 [26] ), .QN(\RegFile/_3895_ ) );
DFF_X1 \RegFile/_8210_ ( .D(\RegFile/_4589_ ), .CK(clock ), .Q(\RegFile/reg_10 [27] ), .QN(\RegFile/_3894_ ) );
DFF_X1 \RegFile/_8211_ ( .D(\RegFile/_4590_ ), .CK(clock ), .Q(\RegFile/reg_10 [28] ), .QN(\RegFile/_3893_ ) );
DFF_X1 \RegFile/_8212_ ( .D(\RegFile/_4591_ ), .CK(clock ), .Q(\RegFile/reg_10 [29] ), .QN(\RegFile/_3892_ ) );
DFF_X1 \RegFile/_8213_ ( .D(\RegFile/_4592_ ), .CK(clock ), .Q(\RegFile/reg_10 [30] ), .QN(\RegFile/_3891_ ) );
DFF_X1 \RegFile/_8214_ ( .D(\RegFile/_4593_ ), .CK(clock ), .Q(\RegFile/reg_10 [31] ), .QN(\RegFile/_3890_ ) );
DFF_X1 \RegFile/_8215_ ( .D(\RegFile/_4594_ ), .CK(clock ), .Q(\RegFile/reg_11 [0] ), .QN(\RegFile/_3889_ ) );
DFF_X1 \RegFile/_8216_ ( .D(\RegFile/_4595_ ), .CK(clock ), .Q(\RegFile/reg_11 [1] ), .QN(\RegFile/_3888_ ) );
DFF_X1 \RegFile/_8217_ ( .D(\RegFile/_4596_ ), .CK(clock ), .Q(\RegFile/reg_11 [2] ), .QN(\RegFile/_3887_ ) );
DFF_X1 \RegFile/_8218_ ( .D(\RegFile/_4597_ ), .CK(clock ), .Q(\RegFile/reg_11 [3] ), .QN(\RegFile/_3886_ ) );
DFF_X1 \RegFile/_8219_ ( .D(\RegFile/_4598_ ), .CK(clock ), .Q(\RegFile/reg_11 [4] ), .QN(\RegFile/_3885_ ) );
DFF_X1 \RegFile/_8220_ ( .D(\RegFile/_4599_ ), .CK(clock ), .Q(\RegFile/reg_11 [5] ), .QN(\RegFile/_3884_ ) );
DFF_X1 \RegFile/_8221_ ( .D(\RegFile/_4600_ ), .CK(clock ), .Q(\RegFile/reg_11 [6] ), .QN(\RegFile/_3883_ ) );
DFF_X1 \RegFile/_8222_ ( .D(\RegFile/_4601_ ), .CK(clock ), .Q(\RegFile/reg_11 [7] ), .QN(\RegFile/_3882_ ) );
DFF_X1 \RegFile/_8223_ ( .D(\RegFile/_4602_ ), .CK(clock ), .Q(\RegFile/reg_11 [8] ), .QN(\RegFile/_3881_ ) );
DFF_X1 \RegFile/_8224_ ( .D(\RegFile/_4603_ ), .CK(clock ), .Q(\RegFile/reg_11 [9] ), .QN(\RegFile/_3880_ ) );
DFF_X1 \RegFile/_8225_ ( .D(\RegFile/_4604_ ), .CK(clock ), .Q(\RegFile/reg_11 [10] ), .QN(\RegFile/_3879_ ) );
DFF_X1 \RegFile/_8226_ ( .D(\RegFile/_4605_ ), .CK(clock ), .Q(\RegFile/reg_11 [11] ), .QN(\RegFile/_3878_ ) );
DFF_X1 \RegFile/_8227_ ( .D(\RegFile/_4606_ ), .CK(clock ), .Q(\RegFile/reg_11 [12] ), .QN(\RegFile/_3877_ ) );
DFF_X1 \RegFile/_8228_ ( .D(\RegFile/_4607_ ), .CK(clock ), .Q(\RegFile/reg_11 [13] ), .QN(\RegFile/_3876_ ) );
DFF_X1 \RegFile/_8229_ ( .D(\RegFile/_4608_ ), .CK(clock ), .Q(\RegFile/reg_11 [14] ), .QN(\RegFile/_3875_ ) );
DFF_X1 \RegFile/_8230_ ( .D(\RegFile/_4609_ ), .CK(clock ), .Q(\RegFile/reg_11 [15] ), .QN(\RegFile/_3874_ ) );
DFF_X1 \RegFile/_8231_ ( .D(\RegFile/_4610_ ), .CK(clock ), .Q(\RegFile/reg_11 [16] ), .QN(\RegFile/_3873_ ) );
DFF_X1 \RegFile/_8232_ ( .D(\RegFile/_4611_ ), .CK(clock ), .Q(\RegFile/reg_11 [17] ), .QN(\RegFile/_3872_ ) );
DFF_X1 \RegFile/_8233_ ( .D(\RegFile/_4612_ ), .CK(clock ), .Q(\RegFile/reg_11 [18] ), .QN(\RegFile/_3871_ ) );
DFF_X1 \RegFile/_8234_ ( .D(\RegFile/_4613_ ), .CK(clock ), .Q(\RegFile/reg_11 [19] ), .QN(\RegFile/_3870_ ) );
DFF_X1 \RegFile/_8235_ ( .D(\RegFile/_4614_ ), .CK(clock ), .Q(\RegFile/reg_11 [20] ), .QN(\RegFile/_3869_ ) );
DFF_X1 \RegFile/_8236_ ( .D(\RegFile/_4615_ ), .CK(clock ), .Q(\RegFile/reg_11 [21] ), .QN(\RegFile/_3868_ ) );
DFF_X1 \RegFile/_8237_ ( .D(\RegFile/_4616_ ), .CK(clock ), .Q(\RegFile/reg_11 [22] ), .QN(\RegFile/_3867_ ) );
DFF_X1 \RegFile/_8238_ ( .D(\RegFile/_4617_ ), .CK(clock ), .Q(\RegFile/reg_11 [23] ), .QN(\RegFile/_3866_ ) );
DFF_X1 \RegFile/_8239_ ( .D(\RegFile/_4618_ ), .CK(clock ), .Q(\RegFile/reg_11 [24] ), .QN(\RegFile/_3865_ ) );
DFF_X1 \RegFile/_8240_ ( .D(\RegFile/_4619_ ), .CK(clock ), .Q(\RegFile/reg_11 [25] ), .QN(\RegFile/_3864_ ) );
DFF_X1 \RegFile/_8241_ ( .D(\RegFile/_4620_ ), .CK(clock ), .Q(\RegFile/reg_11 [26] ), .QN(\RegFile/_3863_ ) );
DFF_X1 \RegFile/_8242_ ( .D(\RegFile/_4621_ ), .CK(clock ), .Q(\RegFile/reg_11 [27] ), .QN(\RegFile/_3862_ ) );
DFF_X1 \RegFile/_8243_ ( .D(\RegFile/_4622_ ), .CK(clock ), .Q(\RegFile/reg_11 [28] ), .QN(\RegFile/_3861_ ) );
DFF_X1 \RegFile/_8244_ ( .D(\RegFile/_4623_ ), .CK(clock ), .Q(\RegFile/reg_11 [29] ), .QN(\RegFile/_3860_ ) );
DFF_X1 \RegFile/_8245_ ( .D(\RegFile/_4624_ ), .CK(clock ), .Q(\RegFile/reg_11 [30] ), .QN(\RegFile/_3859_ ) );
DFF_X1 \RegFile/_8246_ ( .D(\RegFile/_4625_ ), .CK(clock ), .Q(\RegFile/reg_11 [31] ), .QN(\RegFile/_3858_ ) );
DFF_X1 \RegFile/_8247_ ( .D(\RegFile/_4626_ ), .CK(clock ), .Q(\RegFile/reg_12 [0] ), .QN(\RegFile/_3857_ ) );
DFF_X1 \RegFile/_8248_ ( .D(\RegFile/_4627_ ), .CK(clock ), .Q(\RegFile/reg_12 [1] ), .QN(\RegFile/_3856_ ) );
DFF_X1 \RegFile/_8249_ ( .D(\RegFile/_4628_ ), .CK(clock ), .Q(\RegFile/reg_12 [2] ), .QN(\RegFile/_3855_ ) );
DFF_X1 \RegFile/_8250_ ( .D(\RegFile/_4629_ ), .CK(clock ), .Q(\RegFile/reg_12 [3] ), .QN(\RegFile/_3854_ ) );
DFF_X1 \RegFile/_8251_ ( .D(\RegFile/_4630_ ), .CK(clock ), .Q(\RegFile/reg_12 [4] ), .QN(\RegFile/_3853_ ) );
DFF_X1 \RegFile/_8252_ ( .D(\RegFile/_4631_ ), .CK(clock ), .Q(\RegFile/reg_12 [5] ), .QN(\RegFile/_3852_ ) );
DFF_X1 \RegFile/_8253_ ( .D(\RegFile/_4632_ ), .CK(clock ), .Q(\RegFile/reg_12 [6] ), .QN(\RegFile/_3851_ ) );
DFF_X1 \RegFile/_8254_ ( .D(\RegFile/_4633_ ), .CK(clock ), .Q(\RegFile/reg_12 [7] ), .QN(\RegFile/_3850_ ) );
DFF_X1 \RegFile/_8255_ ( .D(\RegFile/_4634_ ), .CK(clock ), .Q(\RegFile/reg_12 [8] ), .QN(\RegFile/_3849_ ) );
DFF_X1 \RegFile/_8256_ ( .D(\RegFile/_4635_ ), .CK(clock ), .Q(\RegFile/reg_12 [9] ), .QN(\RegFile/_3848_ ) );
DFF_X1 \RegFile/_8257_ ( .D(\RegFile/_4636_ ), .CK(clock ), .Q(\RegFile/reg_12 [10] ), .QN(\RegFile/_3847_ ) );
DFF_X1 \RegFile/_8258_ ( .D(\RegFile/_4637_ ), .CK(clock ), .Q(\RegFile/reg_12 [11] ), .QN(\RegFile/_3846_ ) );
DFF_X1 \RegFile/_8259_ ( .D(\RegFile/_4638_ ), .CK(clock ), .Q(\RegFile/reg_12 [12] ), .QN(\RegFile/_3845_ ) );
DFF_X1 \RegFile/_8260_ ( .D(\RegFile/_4639_ ), .CK(clock ), .Q(\RegFile/reg_12 [13] ), .QN(\RegFile/_3844_ ) );
DFF_X1 \RegFile/_8261_ ( .D(\RegFile/_4640_ ), .CK(clock ), .Q(\RegFile/reg_12 [14] ), .QN(\RegFile/_3843_ ) );
DFF_X1 \RegFile/_8262_ ( .D(\RegFile/_4641_ ), .CK(clock ), .Q(\RegFile/reg_12 [15] ), .QN(\RegFile/_3842_ ) );
DFF_X1 \RegFile/_8263_ ( .D(\RegFile/_4642_ ), .CK(clock ), .Q(\RegFile/reg_12 [16] ), .QN(\RegFile/_3841_ ) );
DFF_X1 \RegFile/_8264_ ( .D(\RegFile/_4643_ ), .CK(clock ), .Q(\RegFile/reg_12 [17] ), .QN(\RegFile/_3840_ ) );
DFF_X1 \RegFile/_8265_ ( .D(\RegFile/_4644_ ), .CK(clock ), .Q(\RegFile/reg_12 [18] ), .QN(\RegFile/_3839_ ) );
DFF_X1 \RegFile/_8266_ ( .D(\RegFile/_4645_ ), .CK(clock ), .Q(\RegFile/reg_12 [19] ), .QN(\RegFile/_3838_ ) );
DFF_X1 \RegFile/_8267_ ( .D(\RegFile/_4646_ ), .CK(clock ), .Q(\RegFile/reg_12 [20] ), .QN(\RegFile/_3837_ ) );
DFF_X1 \RegFile/_8268_ ( .D(\RegFile/_4647_ ), .CK(clock ), .Q(\RegFile/reg_12 [21] ), .QN(\RegFile/_3836_ ) );
DFF_X1 \RegFile/_8269_ ( .D(\RegFile/_4648_ ), .CK(clock ), .Q(\RegFile/reg_12 [22] ), .QN(\RegFile/_3835_ ) );
DFF_X1 \RegFile/_8270_ ( .D(\RegFile/_4649_ ), .CK(clock ), .Q(\RegFile/reg_12 [23] ), .QN(\RegFile/_3834_ ) );
DFF_X1 \RegFile/_8271_ ( .D(\RegFile/_4650_ ), .CK(clock ), .Q(\RegFile/reg_12 [24] ), .QN(\RegFile/_3833_ ) );
DFF_X1 \RegFile/_8272_ ( .D(\RegFile/_4651_ ), .CK(clock ), .Q(\RegFile/reg_12 [25] ), .QN(\RegFile/_3832_ ) );
DFF_X1 \RegFile/_8273_ ( .D(\RegFile/_4652_ ), .CK(clock ), .Q(\RegFile/reg_12 [26] ), .QN(\RegFile/_3831_ ) );
DFF_X1 \RegFile/_8274_ ( .D(\RegFile/_4653_ ), .CK(clock ), .Q(\RegFile/reg_12 [27] ), .QN(\RegFile/_3830_ ) );
DFF_X1 \RegFile/_8275_ ( .D(\RegFile/_4654_ ), .CK(clock ), .Q(\RegFile/reg_12 [28] ), .QN(\RegFile/_3829_ ) );
DFF_X1 \RegFile/_8276_ ( .D(\RegFile/_4655_ ), .CK(clock ), .Q(\RegFile/reg_12 [29] ), .QN(\RegFile/_3828_ ) );
DFF_X1 \RegFile/_8277_ ( .D(\RegFile/_4656_ ), .CK(clock ), .Q(\RegFile/reg_12 [30] ), .QN(\RegFile/_3827_ ) );
DFF_X1 \RegFile/_8278_ ( .D(\RegFile/_4657_ ), .CK(clock ), .Q(\RegFile/reg_12 [31] ), .QN(\RegFile/_3826_ ) );
DFF_X1 \RegFile/_8279_ ( .D(\RegFile/_4658_ ), .CK(clock ), .Q(\RegFile/reg_13 [0] ), .QN(\RegFile/_3825_ ) );
DFF_X1 \RegFile/_8280_ ( .D(\RegFile/_4659_ ), .CK(clock ), .Q(\RegFile/reg_13 [1] ), .QN(\RegFile/_3824_ ) );
DFF_X1 \RegFile/_8281_ ( .D(\RegFile/_4660_ ), .CK(clock ), .Q(\RegFile/reg_13 [2] ), .QN(\RegFile/_3823_ ) );
DFF_X1 \RegFile/_8282_ ( .D(\RegFile/_4661_ ), .CK(clock ), .Q(\RegFile/reg_13 [3] ), .QN(\RegFile/_3822_ ) );
DFF_X1 \RegFile/_8283_ ( .D(\RegFile/_4662_ ), .CK(clock ), .Q(\RegFile/reg_13 [4] ), .QN(\RegFile/_3821_ ) );
DFF_X1 \RegFile/_8284_ ( .D(\RegFile/_4663_ ), .CK(clock ), .Q(\RegFile/reg_13 [5] ), .QN(\RegFile/_3820_ ) );
DFF_X1 \RegFile/_8285_ ( .D(\RegFile/_4664_ ), .CK(clock ), .Q(\RegFile/reg_13 [6] ), .QN(\RegFile/_3819_ ) );
DFF_X1 \RegFile/_8286_ ( .D(\RegFile/_4665_ ), .CK(clock ), .Q(\RegFile/reg_13 [7] ), .QN(\RegFile/_3818_ ) );
DFF_X1 \RegFile/_8287_ ( .D(\RegFile/_4666_ ), .CK(clock ), .Q(\RegFile/reg_13 [8] ), .QN(\RegFile/_3817_ ) );
DFF_X1 \RegFile/_8288_ ( .D(\RegFile/_4667_ ), .CK(clock ), .Q(\RegFile/reg_13 [9] ), .QN(\RegFile/_3816_ ) );
DFF_X1 \RegFile/_8289_ ( .D(\RegFile/_4668_ ), .CK(clock ), .Q(\RegFile/reg_13 [10] ), .QN(\RegFile/_3815_ ) );
DFF_X1 \RegFile/_8290_ ( .D(\RegFile/_4669_ ), .CK(clock ), .Q(\RegFile/reg_13 [11] ), .QN(\RegFile/_3814_ ) );
DFF_X1 \RegFile/_8291_ ( .D(\RegFile/_4670_ ), .CK(clock ), .Q(\RegFile/reg_13 [12] ), .QN(\RegFile/_3813_ ) );
DFF_X1 \RegFile/_8292_ ( .D(\RegFile/_4671_ ), .CK(clock ), .Q(\RegFile/reg_13 [13] ), .QN(\RegFile/_3812_ ) );
DFF_X1 \RegFile/_8293_ ( .D(\RegFile/_4672_ ), .CK(clock ), .Q(\RegFile/reg_13 [14] ), .QN(\RegFile/_3811_ ) );
DFF_X1 \RegFile/_8294_ ( .D(\RegFile/_4673_ ), .CK(clock ), .Q(\RegFile/reg_13 [15] ), .QN(\RegFile/_3810_ ) );
DFF_X1 \RegFile/_8295_ ( .D(\RegFile/_4674_ ), .CK(clock ), .Q(\RegFile/reg_13 [16] ), .QN(\RegFile/_3809_ ) );
DFF_X1 \RegFile/_8296_ ( .D(\RegFile/_4675_ ), .CK(clock ), .Q(\RegFile/reg_13 [17] ), .QN(\RegFile/_3808_ ) );
DFF_X1 \RegFile/_8297_ ( .D(\RegFile/_4676_ ), .CK(clock ), .Q(\RegFile/reg_13 [18] ), .QN(\RegFile/_3807_ ) );
DFF_X1 \RegFile/_8298_ ( .D(\RegFile/_4677_ ), .CK(clock ), .Q(\RegFile/reg_13 [19] ), .QN(\RegFile/_3806_ ) );
DFF_X1 \RegFile/_8299_ ( .D(\RegFile/_4678_ ), .CK(clock ), .Q(\RegFile/reg_13 [20] ), .QN(\RegFile/_3805_ ) );
DFF_X1 \RegFile/_8300_ ( .D(\RegFile/_4679_ ), .CK(clock ), .Q(\RegFile/reg_13 [21] ), .QN(\RegFile/_3804_ ) );
DFF_X1 \RegFile/_8301_ ( .D(\RegFile/_4680_ ), .CK(clock ), .Q(\RegFile/reg_13 [22] ), .QN(\RegFile/_3803_ ) );
DFF_X1 \RegFile/_8302_ ( .D(\RegFile/_4681_ ), .CK(clock ), .Q(\RegFile/reg_13 [23] ), .QN(\RegFile/_3802_ ) );
DFF_X1 \RegFile/_8303_ ( .D(\RegFile/_4682_ ), .CK(clock ), .Q(\RegFile/reg_13 [24] ), .QN(\RegFile/_3801_ ) );
DFF_X1 \RegFile/_8304_ ( .D(\RegFile/_4683_ ), .CK(clock ), .Q(\RegFile/reg_13 [25] ), .QN(\RegFile/_3800_ ) );
DFF_X1 \RegFile/_8305_ ( .D(\RegFile/_4684_ ), .CK(clock ), .Q(\RegFile/reg_13 [26] ), .QN(\RegFile/_3799_ ) );
DFF_X1 \RegFile/_8306_ ( .D(\RegFile/_4685_ ), .CK(clock ), .Q(\RegFile/reg_13 [27] ), .QN(\RegFile/_3798_ ) );
DFF_X1 \RegFile/_8307_ ( .D(\RegFile/_4686_ ), .CK(clock ), .Q(\RegFile/reg_13 [28] ), .QN(\RegFile/_3797_ ) );
DFF_X1 \RegFile/_8308_ ( .D(\RegFile/_4687_ ), .CK(clock ), .Q(\RegFile/reg_13 [29] ), .QN(\RegFile/_3796_ ) );
DFF_X1 \RegFile/_8309_ ( .D(\RegFile/_4688_ ), .CK(clock ), .Q(\RegFile/reg_13 [30] ), .QN(\RegFile/_3795_ ) );
DFF_X1 \RegFile/_8310_ ( .D(\RegFile/_4689_ ), .CK(clock ), .Q(\RegFile/reg_13 [31] ), .QN(\RegFile/_3794_ ) );
DFF_X1 \RegFile/_8311_ ( .D(\RegFile/_4690_ ), .CK(clock ), .Q(\RegFile/reg_14 [0] ), .QN(\RegFile/_0047_ ) );
DFF_X1 \RegFile/_8312_ ( .D(\RegFile/_4691_ ), .CK(clock ), .Q(\RegFile/reg_14 [1] ), .QN(\RegFile/_0049_ ) );
DFF_X1 \RegFile/_8313_ ( .D(\RegFile/_4692_ ), .CK(clock ), .Q(\RegFile/reg_14 [2] ), .QN(\RegFile/_0051_ ) );
DFF_X1 \RegFile/_8314_ ( .D(\RegFile/_4693_ ), .CK(clock ), .Q(\RegFile/reg_14 [3] ), .QN(\RegFile/_0053_ ) );
DFF_X1 \RegFile/_8315_ ( .D(\RegFile/_4694_ ), .CK(clock ), .Q(\RegFile/reg_14 [4] ), .QN(\RegFile/_0055_ ) );
DFF_X1 \RegFile/_8316_ ( .D(\RegFile/_4695_ ), .CK(clock ), .Q(\RegFile/reg_14 [5] ), .QN(\RegFile/_0057_ ) );
DFF_X1 \RegFile/_8317_ ( .D(\RegFile/_4696_ ), .CK(clock ), .Q(\RegFile/reg_14 [6] ), .QN(\RegFile/_0059_ ) );
DFF_X1 \RegFile/_8318_ ( .D(\RegFile/_4697_ ), .CK(clock ), .Q(\RegFile/reg_14 [7] ), .QN(\RegFile/_0061_ ) );
DFF_X1 \RegFile/_8319_ ( .D(\RegFile/_4698_ ), .CK(clock ), .Q(\RegFile/reg_14 [8] ), .QN(\RegFile/_0063_ ) );
DFF_X1 \RegFile/_8320_ ( .D(\RegFile/_4699_ ), .CK(clock ), .Q(\RegFile/reg_14 [9] ), .QN(\RegFile/_0001_ ) );
DFF_X1 \RegFile/_8321_ ( .D(\RegFile/_4700_ ), .CK(clock ), .Q(\RegFile/reg_14 [10] ), .QN(\RegFile/_0003_ ) );
DFF_X1 \RegFile/_8322_ ( .D(\RegFile/_4701_ ), .CK(clock ), .Q(\RegFile/reg_14 [11] ), .QN(\RegFile/_0005_ ) );
DFF_X1 \RegFile/_8323_ ( .D(\RegFile/_4702_ ), .CK(clock ), .Q(\RegFile/reg_14 [12] ), .QN(\RegFile/_0007_ ) );
DFF_X1 \RegFile/_8324_ ( .D(\RegFile/_4703_ ), .CK(clock ), .Q(\RegFile/reg_14 [13] ), .QN(\RegFile/_0009_ ) );
DFF_X1 \RegFile/_8325_ ( .D(\RegFile/_4704_ ), .CK(clock ), .Q(\RegFile/reg_14 [14] ), .QN(\RegFile/_0011_ ) );
DFF_X1 \RegFile/_8326_ ( .D(\RegFile/_4705_ ), .CK(clock ), .Q(\RegFile/reg_14 [15] ), .QN(\RegFile/_0013_ ) );
DFF_X1 \RegFile/_8327_ ( .D(\RegFile/_4706_ ), .CK(clock ), .Q(\RegFile/reg_14 [16] ), .QN(\RegFile/_0015_ ) );
DFF_X1 \RegFile/_8328_ ( .D(\RegFile/_4707_ ), .CK(clock ), .Q(\RegFile/reg_14 [17] ), .QN(\RegFile/_0017_ ) );
DFF_X1 \RegFile/_8329_ ( .D(\RegFile/_4708_ ), .CK(clock ), .Q(\RegFile/reg_14 [18] ), .QN(\RegFile/_0019_ ) );
DFF_X1 \RegFile/_8330_ ( .D(\RegFile/_4709_ ), .CK(clock ), .Q(\RegFile/reg_14 [19] ), .QN(\RegFile/_0021_ ) );
DFF_X1 \RegFile/_8331_ ( .D(\RegFile/_4710_ ), .CK(clock ), .Q(\RegFile/reg_14 [20] ), .QN(\RegFile/_0023_ ) );
DFF_X1 \RegFile/_8332_ ( .D(\RegFile/_4711_ ), .CK(clock ), .Q(\RegFile/reg_14 [21] ), .QN(\RegFile/_0025_ ) );
DFF_X1 \RegFile/_8333_ ( .D(\RegFile/_4712_ ), .CK(clock ), .Q(\RegFile/reg_14 [22] ), .QN(\RegFile/_0027_ ) );
DFF_X1 \RegFile/_8334_ ( .D(\RegFile/_4713_ ), .CK(clock ), .Q(\RegFile/reg_14 [23] ), .QN(\RegFile/_0029_ ) );
DFF_X1 \RegFile/_8335_ ( .D(\RegFile/_4714_ ), .CK(clock ), .Q(\RegFile/reg_14 [24] ), .QN(\RegFile/_0031_ ) );
DFF_X1 \RegFile/_8336_ ( .D(\RegFile/_4715_ ), .CK(clock ), .Q(\RegFile/reg_14 [25] ), .QN(\RegFile/_0033_ ) );
DFF_X1 \RegFile/_8337_ ( .D(\RegFile/_4716_ ), .CK(clock ), .Q(\RegFile/reg_14 [26] ), .QN(\RegFile/_0035_ ) );
DFF_X1 \RegFile/_8338_ ( .D(\RegFile/_4717_ ), .CK(clock ), .Q(\RegFile/reg_14 [27] ), .QN(\RegFile/_0037_ ) );
DFF_X1 \RegFile/_8339_ ( .D(\RegFile/_4718_ ), .CK(clock ), .Q(\RegFile/reg_14 [28] ), .QN(\RegFile/_0039_ ) );
DFF_X1 \RegFile/_8340_ ( .D(\RegFile/_4719_ ), .CK(clock ), .Q(\RegFile/reg_14 [29] ), .QN(\RegFile/_0041_ ) );
DFF_X1 \RegFile/_8341_ ( .D(\RegFile/_4720_ ), .CK(clock ), .Q(\RegFile/reg_14 [30] ), .QN(\RegFile/_0043_ ) );
DFF_X1 \RegFile/_8342_ ( .D(\RegFile/_4721_ ), .CK(clock ), .Q(\RegFile/reg_14 [31] ), .QN(\RegFile/_0045_ ) );
DFF_X1 \RegFile/_8343_ ( .D(\RegFile/_4722_ ), .CK(clock ), .Q(\RegFile/reg_15 [0] ), .QN(\RegFile/_0046_ ) );
DFF_X1 \RegFile/_8344_ ( .D(\RegFile/_4723_ ), .CK(clock ), .Q(\RegFile/reg_15 [1] ), .QN(\RegFile/_0048_ ) );
DFF_X1 \RegFile/_8345_ ( .D(\RegFile/_4724_ ), .CK(clock ), .Q(\RegFile/reg_15 [2] ), .QN(\RegFile/_0050_ ) );
DFF_X1 \RegFile/_8346_ ( .D(\RegFile/_4725_ ), .CK(clock ), .Q(\RegFile/reg_15 [3] ), .QN(\RegFile/_0052_ ) );
DFF_X1 \RegFile/_8347_ ( .D(\RegFile/_4726_ ), .CK(clock ), .Q(\RegFile/reg_15 [4] ), .QN(\RegFile/_0054_ ) );
DFF_X1 \RegFile/_8348_ ( .D(\RegFile/_4727_ ), .CK(clock ), .Q(\RegFile/reg_15 [5] ), .QN(\RegFile/_0056_ ) );
DFF_X1 \RegFile/_8349_ ( .D(\RegFile/_4728_ ), .CK(clock ), .Q(\RegFile/reg_15 [6] ), .QN(\RegFile/_0058_ ) );
DFF_X1 \RegFile/_8350_ ( .D(\RegFile/_4729_ ), .CK(clock ), .Q(\RegFile/reg_15 [7] ), .QN(\RegFile/_0060_ ) );
DFF_X1 \RegFile/_8351_ ( .D(\RegFile/_4730_ ), .CK(clock ), .Q(\RegFile/reg_15 [8] ), .QN(\RegFile/_0062_ ) );
DFF_X1 \RegFile/_8352_ ( .D(\RegFile/_4731_ ), .CK(clock ), .Q(\RegFile/reg_15 [9] ), .QN(\RegFile/_0000_ ) );
DFF_X1 \RegFile/_8353_ ( .D(\RegFile/_4732_ ), .CK(clock ), .Q(\RegFile/reg_15 [10] ), .QN(\RegFile/_0002_ ) );
DFF_X1 \RegFile/_8354_ ( .D(\RegFile/_4733_ ), .CK(clock ), .Q(\RegFile/reg_15 [11] ), .QN(\RegFile/_0004_ ) );
DFF_X1 \RegFile/_8355_ ( .D(\RegFile/_4734_ ), .CK(clock ), .Q(\RegFile/reg_15 [12] ), .QN(\RegFile/_0006_ ) );
DFF_X1 \RegFile/_8356_ ( .D(\RegFile/_4735_ ), .CK(clock ), .Q(\RegFile/reg_15 [13] ), .QN(\RegFile/_0008_ ) );
DFF_X1 \RegFile/_8357_ ( .D(\RegFile/_4736_ ), .CK(clock ), .Q(\RegFile/reg_15 [14] ), .QN(\RegFile/_0010_ ) );
DFF_X1 \RegFile/_8358_ ( .D(\RegFile/_4737_ ), .CK(clock ), .Q(\RegFile/reg_15 [15] ), .QN(\RegFile/_0012_ ) );
DFF_X1 \RegFile/_8359_ ( .D(\RegFile/_4738_ ), .CK(clock ), .Q(\RegFile/reg_15 [16] ), .QN(\RegFile/_0014_ ) );
DFF_X1 \RegFile/_8360_ ( .D(\RegFile/_4739_ ), .CK(clock ), .Q(\RegFile/reg_15 [17] ), .QN(\RegFile/_0016_ ) );
DFF_X1 \RegFile/_8361_ ( .D(\RegFile/_4740_ ), .CK(clock ), .Q(\RegFile/reg_15 [18] ), .QN(\RegFile/_0018_ ) );
DFF_X1 \RegFile/_8362_ ( .D(\RegFile/_4741_ ), .CK(clock ), .Q(\RegFile/reg_15 [19] ), .QN(\RegFile/_0020_ ) );
DFF_X1 \RegFile/_8363_ ( .D(\RegFile/_4742_ ), .CK(clock ), .Q(\RegFile/reg_15 [20] ), .QN(\RegFile/_0022_ ) );
DFF_X1 \RegFile/_8364_ ( .D(\RegFile/_4743_ ), .CK(clock ), .Q(\RegFile/reg_15 [21] ), .QN(\RegFile/_0024_ ) );
DFF_X1 \RegFile/_8365_ ( .D(\RegFile/_4744_ ), .CK(clock ), .Q(\RegFile/reg_15 [22] ), .QN(\RegFile/_0026_ ) );
DFF_X1 \RegFile/_8366_ ( .D(\RegFile/_4745_ ), .CK(clock ), .Q(\RegFile/reg_15 [23] ), .QN(\RegFile/_0028_ ) );
DFF_X1 \RegFile/_8367_ ( .D(\RegFile/_4746_ ), .CK(clock ), .Q(\RegFile/reg_15 [24] ), .QN(\RegFile/_0030_ ) );
DFF_X1 \RegFile/_8368_ ( .D(\RegFile/_4747_ ), .CK(clock ), .Q(\RegFile/reg_15 [25] ), .QN(\RegFile/_0032_ ) );
DFF_X1 \RegFile/_8369_ ( .D(\RegFile/_4748_ ), .CK(clock ), .Q(\RegFile/reg_15 [26] ), .QN(\RegFile/_0034_ ) );
DFF_X1 \RegFile/_8370_ ( .D(\RegFile/_4749_ ), .CK(clock ), .Q(\RegFile/reg_15 [27] ), .QN(\RegFile/_0036_ ) );
DFF_X1 \RegFile/_8371_ ( .D(\RegFile/_4750_ ), .CK(clock ), .Q(\RegFile/reg_15 [28] ), .QN(\RegFile/_0038_ ) );
DFF_X1 \RegFile/_8372_ ( .D(\RegFile/_4751_ ), .CK(clock ), .Q(\RegFile/reg_15 [29] ), .QN(\RegFile/_0040_ ) );
DFF_X1 \RegFile/_8373_ ( .D(\RegFile/_4752_ ), .CK(clock ), .Q(\RegFile/reg_15 [30] ), .QN(\RegFile/_0042_ ) );
DFF_X1 \RegFile/_8374_ ( .D(\RegFile/_4753_ ), .CK(clock ), .Q(\RegFile/reg_15 [31] ), .QN(\RegFile/_0044_ ) );
BUF_X1 \RegFile/_8375_ ( .A(\_WBU_io_RegFileAccess_wa [1] ), .Z(\RegFile/_0713_ ) );
BUF_X1 \RegFile/_8376_ ( .A(\_WBU_io_RegFileAccess_wa [0] ), .Z(\RegFile/_0712_ ) );
BUF_X1 \RegFile/_8377_ ( .A(\_WBU_io_RegFileAccess_wa [3] ), .Z(\RegFile/_0715_ ) );
BUF_X1 \RegFile/_8378_ ( .A(\_WBU_io_RegFileAccess_wa [2] ), .Z(\RegFile/_0714_ ) );
BUF_X1 \RegFile/_8379_ ( .A(\_IDU_io_RegFileAccess_ra1 [1] ), .Z(\RegFile/_0641_ ) );
BUF_X1 \RegFile/_8380_ ( .A(\_IDU_io_RegFileAccess_ra1 [0] ), .Z(\RegFile/_0640_ ) );
BUF_X1 \RegFile/_8381_ ( .A(\_IDU_io_RegFileAccess_ra1 [3] ), .Z(\RegFile/_0643_ ) );
BUF_X1 \RegFile/_8382_ ( .A(\_IDU_io_RegFileAccess_ra1 [2] ), .Z(\RegFile/_0642_ ) );
BUF_X1 \RegFile/_8383_ ( .A(\RegFile/_0047_ ), .Z(\RegFile/_0111_ ) );
BUF_X1 \RegFile/_8384_ ( .A(\RegFile/reg_13 [0] ), .Z(\RegFile/_3410_ ) );
BUF_X1 \RegFile/_8385_ ( .A(\RegFile/reg_12 [0] ), .Z(\RegFile/_3378_ ) );
BUF_X1 \RegFile/_8386_ ( .A(\RegFile/reg_11 [0] ), .Z(\RegFile/_3346_ ) );
BUF_X1 \RegFile/_8387_ ( .A(\RegFile/reg_10 [0] ), .Z(\RegFile/_3314_ ) );
BUF_X1 \RegFile/_8388_ ( .A(\RegFile/reg_9 [0] ), .Z(\RegFile/_3762_ ) );
BUF_X1 \RegFile/_8389_ ( .A(\RegFile/reg_8 [0] ), .Z(\RegFile/_3730_ ) );
BUF_X1 \RegFile/_8390_ ( .A(\RegFile/reg_7 [0] ), .Z(\RegFile/_3698_ ) );
BUF_X1 \RegFile/_8391_ ( .A(\RegFile/reg_6 [0] ), .Z(\RegFile/_3666_ ) );
BUF_X1 \RegFile/_8392_ ( .A(\RegFile/reg_5 [0] ), .Z(\RegFile/_3634_ ) );
BUF_X1 \RegFile/_8393_ ( .A(\RegFile/reg_4 [0] ), .Z(\RegFile/_3602_ ) );
BUF_X1 \RegFile/_8394_ ( .A(\RegFile/reg_3 [0] ), .Z(\RegFile/_3570_ ) );
BUF_X1 \RegFile/_8395_ ( .A(\RegFile/reg_2 [0] ), .Z(\RegFile/_3538_ ) );
BUF_X1 \RegFile/_8396_ ( .A(\RegFile/reg_1 [0] ), .Z(\RegFile/_3506_ ) );
BUF_X1 \RegFile/_8397_ ( .A(\RegFile/reg_0 [0] ), .Z(\RegFile/_3282_ ) );
BUF_X1 \RegFile/_8398_ ( .A(\RegFile/_0046_ ), .Z(\RegFile/_0110_ ) );
BUF_X1 \RegFile/_8399_ ( .A(\RegFile/_0648_ ), .Z(\_RegFile_io_rd1 [0] ) );
BUF_X1 \RegFile/_8400_ ( .A(\RegFile/_0049_ ), .Z(\RegFile/_0113_ ) );
BUF_X1 \RegFile/_8401_ ( .A(\RegFile/reg_13 [1] ), .Z(\RegFile/_3421_ ) );
BUF_X1 \RegFile/_8402_ ( .A(\RegFile/reg_12 [1] ), .Z(\RegFile/_3389_ ) );
BUF_X1 \RegFile/_8403_ ( .A(\RegFile/reg_11 [1] ), .Z(\RegFile/_3357_ ) );
BUF_X1 \RegFile/_8404_ ( .A(\RegFile/reg_10 [1] ), .Z(\RegFile/_3325_ ) );
BUF_X1 \RegFile/_8405_ ( .A(\RegFile/reg_9 [1] ), .Z(\RegFile/_3773_ ) );
BUF_X1 \RegFile/_8406_ ( .A(\RegFile/reg_8 [1] ), .Z(\RegFile/_3741_ ) );
BUF_X1 \RegFile/_8407_ ( .A(\RegFile/reg_7 [1] ), .Z(\RegFile/_3709_ ) );
BUF_X1 \RegFile/_8408_ ( .A(\RegFile/reg_6 [1] ), .Z(\RegFile/_3677_ ) );
BUF_X1 \RegFile/_8409_ ( .A(\RegFile/reg_5 [1] ), .Z(\RegFile/_3645_ ) );
BUF_X1 \RegFile/_8410_ ( .A(\RegFile/reg_4 [1] ), .Z(\RegFile/_3613_ ) );
BUF_X1 \RegFile/_8411_ ( .A(\RegFile/reg_3 [1] ), .Z(\RegFile/_3581_ ) );
BUF_X1 \RegFile/_8412_ ( .A(\RegFile/reg_2 [1] ), .Z(\RegFile/_3549_ ) );
BUF_X1 \RegFile/_8413_ ( .A(\RegFile/reg_1 [1] ), .Z(\RegFile/_3517_ ) );
BUF_X1 \RegFile/_8414_ ( .A(\RegFile/reg_0 [1] ), .Z(\RegFile/_3293_ ) );
BUF_X1 \RegFile/_8415_ ( .A(\RegFile/_0048_ ), .Z(\RegFile/_0112_ ) );
BUF_X1 \RegFile/_8416_ ( .A(\RegFile/_0659_ ), .Z(\_RegFile_io_rd1 [1] ) );
BUF_X1 \RegFile/_8417_ ( .A(\RegFile/_0051_ ), .Z(\RegFile/_0115_ ) );
BUF_X1 \RegFile/_8418_ ( .A(\RegFile/reg_13 [2] ), .Z(\RegFile/_3432_ ) );
BUF_X1 \RegFile/_8419_ ( .A(\RegFile/reg_12 [2] ), .Z(\RegFile/_3400_ ) );
BUF_X1 \RegFile/_8420_ ( .A(\RegFile/reg_11 [2] ), .Z(\RegFile/_3368_ ) );
BUF_X1 \RegFile/_8421_ ( .A(\RegFile/reg_10 [2] ), .Z(\RegFile/_3336_ ) );
BUF_X1 \RegFile/_8422_ ( .A(\RegFile/reg_9 [2] ), .Z(\RegFile/_3784_ ) );
BUF_X1 \RegFile/_8423_ ( .A(\RegFile/reg_8 [2] ), .Z(\RegFile/_3752_ ) );
BUF_X1 \RegFile/_8424_ ( .A(\RegFile/reg_7 [2] ), .Z(\RegFile/_3720_ ) );
BUF_X1 \RegFile/_8425_ ( .A(\RegFile/reg_6 [2] ), .Z(\RegFile/_3688_ ) );
BUF_X1 \RegFile/_8426_ ( .A(\RegFile/reg_5 [2] ), .Z(\RegFile/_3656_ ) );
BUF_X1 \RegFile/_8427_ ( .A(\RegFile/reg_4 [2] ), .Z(\RegFile/_3624_ ) );
BUF_X1 \RegFile/_8428_ ( .A(\RegFile/reg_3 [2] ), .Z(\RegFile/_3592_ ) );
BUF_X1 \RegFile/_8429_ ( .A(\RegFile/reg_2 [2] ), .Z(\RegFile/_3560_ ) );
BUF_X1 \RegFile/_8430_ ( .A(\RegFile/reg_1 [2] ), .Z(\RegFile/_3528_ ) );
BUF_X1 \RegFile/_8431_ ( .A(\RegFile/reg_0 [2] ), .Z(\RegFile/_3304_ ) );
BUF_X1 \RegFile/_8432_ ( .A(\RegFile/_0050_ ), .Z(\RegFile/_0114_ ) );
BUF_X1 \RegFile/_8433_ ( .A(\RegFile/_0670_ ), .Z(\_RegFile_io_rd1 [2] ) );
BUF_X1 \RegFile/_8434_ ( .A(\RegFile/_0053_ ), .Z(\RegFile/_0117_ ) );
BUF_X1 \RegFile/_8435_ ( .A(\RegFile/reg_13 [3] ), .Z(\RegFile/_3435_ ) );
BUF_X1 \RegFile/_8436_ ( .A(\RegFile/reg_12 [3] ), .Z(\RegFile/_3403_ ) );
BUF_X1 \RegFile/_8437_ ( .A(\RegFile/reg_11 [3] ), .Z(\RegFile/_3371_ ) );
BUF_X1 \RegFile/_8438_ ( .A(\RegFile/reg_10 [3] ), .Z(\RegFile/_3339_ ) );
BUF_X1 \RegFile/_8439_ ( .A(\RegFile/reg_9 [3] ), .Z(\RegFile/_3787_ ) );
BUF_X1 \RegFile/_8440_ ( .A(\RegFile/reg_8 [3] ), .Z(\RegFile/_3755_ ) );
BUF_X1 \RegFile/_8441_ ( .A(\RegFile/reg_7 [3] ), .Z(\RegFile/_3723_ ) );
BUF_X1 \RegFile/_8442_ ( .A(\RegFile/reg_6 [3] ), .Z(\RegFile/_3691_ ) );
BUF_X1 \RegFile/_8443_ ( .A(\RegFile/reg_5 [3] ), .Z(\RegFile/_3659_ ) );
BUF_X1 \RegFile/_8444_ ( .A(\RegFile/reg_4 [3] ), .Z(\RegFile/_3627_ ) );
BUF_X1 \RegFile/_8445_ ( .A(\RegFile/reg_3 [3] ), .Z(\RegFile/_3595_ ) );
BUF_X1 \RegFile/_8446_ ( .A(\RegFile/reg_2 [3] ), .Z(\RegFile/_3563_ ) );
BUF_X1 \RegFile/_8447_ ( .A(\RegFile/reg_1 [3] ), .Z(\RegFile/_3531_ ) );
BUF_X1 \RegFile/_8448_ ( .A(\RegFile/reg_0 [3] ), .Z(\RegFile/_3307_ ) );
BUF_X1 \RegFile/_8449_ ( .A(\RegFile/_0052_ ), .Z(\RegFile/_0116_ ) );
BUF_X1 \RegFile/_8450_ ( .A(\RegFile/_0673_ ), .Z(\_RegFile_io_rd1 [3] ) );
BUF_X1 \RegFile/_8451_ ( .A(\RegFile/_0055_ ), .Z(\RegFile/_0119_ ) );
BUF_X1 \RegFile/_8452_ ( .A(\RegFile/reg_13 [4] ), .Z(\RegFile/_3436_ ) );
BUF_X1 \RegFile/_8453_ ( .A(\RegFile/reg_12 [4] ), .Z(\RegFile/_3404_ ) );
BUF_X1 \RegFile/_8454_ ( .A(\RegFile/reg_11 [4] ), .Z(\RegFile/_3372_ ) );
BUF_X1 \RegFile/_8455_ ( .A(\RegFile/reg_10 [4] ), .Z(\RegFile/_3340_ ) );
BUF_X1 \RegFile/_8456_ ( .A(\RegFile/reg_9 [4] ), .Z(\RegFile/_3788_ ) );
BUF_X1 \RegFile/_8457_ ( .A(\RegFile/reg_8 [4] ), .Z(\RegFile/_3756_ ) );
BUF_X1 \RegFile/_8458_ ( .A(\RegFile/reg_7 [4] ), .Z(\RegFile/_3724_ ) );
BUF_X1 \RegFile/_8459_ ( .A(\RegFile/reg_6 [4] ), .Z(\RegFile/_3692_ ) );
BUF_X1 \RegFile/_8460_ ( .A(\RegFile/reg_5 [4] ), .Z(\RegFile/_3660_ ) );
BUF_X1 \RegFile/_8461_ ( .A(\RegFile/reg_4 [4] ), .Z(\RegFile/_3628_ ) );
BUF_X1 \RegFile/_8462_ ( .A(\RegFile/reg_3 [4] ), .Z(\RegFile/_3596_ ) );
BUF_X1 \RegFile/_8463_ ( .A(\RegFile/reg_2 [4] ), .Z(\RegFile/_3564_ ) );
BUF_X1 \RegFile/_8464_ ( .A(\RegFile/reg_1 [4] ), .Z(\RegFile/_3532_ ) );
BUF_X1 \RegFile/_8465_ ( .A(\RegFile/reg_0 [4] ), .Z(\RegFile/_3308_ ) );
BUF_X1 \RegFile/_8466_ ( .A(\RegFile/_0054_ ), .Z(\RegFile/_0118_ ) );
BUF_X1 \RegFile/_8467_ ( .A(\RegFile/_0674_ ), .Z(\_RegFile_io_rd1 [4] ) );
BUF_X1 \RegFile/_8468_ ( .A(\RegFile/_0057_ ), .Z(\RegFile/_0121_ ) );
BUF_X1 \RegFile/_8469_ ( .A(\RegFile/reg_13 [5] ), .Z(\RegFile/_3437_ ) );
BUF_X1 \RegFile/_8470_ ( .A(\RegFile/reg_12 [5] ), .Z(\RegFile/_3405_ ) );
BUF_X1 \RegFile/_8471_ ( .A(\RegFile/reg_11 [5] ), .Z(\RegFile/_3373_ ) );
BUF_X1 \RegFile/_8472_ ( .A(\RegFile/reg_10 [5] ), .Z(\RegFile/_3341_ ) );
BUF_X1 \RegFile/_8473_ ( .A(\RegFile/reg_9 [5] ), .Z(\RegFile/_3789_ ) );
BUF_X1 \RegFile/_8474_ ( .A(\RegFile/reg_8 [5] ), .Z(\RegFile/_3757_ ) );
BUF_X1 \RegFile/_8475_ ( .A(\RegFile/reg_7 [5] ), .Z(\RegFile/_3725_ ) );
BUF_X1 \RegFile/_8476_ ( .A(\RegFile/reg_6 [5] ), .Z(\RegFile/_3693_ ) );
BUF_X1 \RegFile/_8477_ ( .A(\RegFile/reg_5 [5] ), .Z(\RegFile/_3661_ ) );
BUF_X1 \RegFile/_8478_ ( .A(\RegFile/reg_4 [5] ), .Z(\RegFile/_3629_ ) );
BUF_X1 \RegFile/_8479_ ( .A(\RegFile/reg_3 [5] ), .Z(\RegFile/_3597_ ) );
BUF_X1 \RegFile/_8480_ ( .A(\RegFile/reg_2 [5] ), .Z(\RegFile/_3565_ ) );
BUF_X1 \RegFile/_8481_ ( .A(\RegFile/reg_1 [5] ), .Z(\RegFile/_3533_ ) );
BUF_X1 \RegFile/_8482_ ( .A(\RegFile/reg_0 [5] ), .Z(\RegFile/_3309_ ) );
BUF_X1 \RegFile/_8483_ ( .A(\RegFile/_0056_ ), .Z(\RegFile/_0120_ ) );
BUF_X1 \RegFile/_8484_ ( .A(\RegFile/_0675_ ), .Z(\_RegFile_io_rd1 [5] ) );
BUF_X1 \RegFile/_8485_ ( .A(\RegFile/_0059_ ), .Z(\RegFile/_0123_ ) );
BUF_X1 \RegFile/_8486_ ( .A(\RegFile/reg_13 [6] ), .Z(\RegFile/_3438_ ) );
BUF_X1 \RegFile/_8487_ ( .A(\RegFile/reg_12 [6] ), .Z(\RegFile/_3406_ ) );
BUF_X1 \RegFile/_8488_ ( .A(\RegFile/reg_11 [6] ), .Z(\RegFile/_3374_ ) );
BUF_X1 \RegFile/_8489_ ( .A(\RegFile/reg_10 [6] ), .Z(\RegFile/_3342_ ) );
BUF_X1 \RegFile/_8490_ ( .A(\RegFile/reg_9 [6] ), .Z(\RegFile/_3790_ ) );
BUF_X1 \RegFile/_8491_ ( .A(\RegFile/reg_8 [6] ), .Z(\RegFile/_3758_ ) );
BUF_X1 \RegFile/_8492_ ( .A(\RegFile/reg_7 [6] ), .Z(\RegFile/_3726_ ) );
BUF_X1 \RegFile/_8493_ ( .A(\RegFile/reg_6 [6] ), .Z(\RegFile/_3694_ ) );
BUF_X1 \RegFile/_8494_ ( .A(\RegFile/reg_5 [6] ), .Z(\RegFile/_3662_ ) );
BUF_X1 \RegFile/_8495_ ( .A(\RegFile/reg_4 [6] ), .Z(\RegFile/_3630_ ) );
BUF_X1 \RegFile/_8496_ ( .A(\RegFile/reg_3 [6] ), .Z(\RegFile/_3598_ ) );
BUF_X1 \RegFile/_8497_ ( .A(\RegFile/reg_2 [6] ), .Z(\RegFile/_3566_ ) );
BUF_X1 \RegFile/_8498_ ( .A(\RegFile/reg_1 [6] ), .Z(\RegFile/_3534_ ) );
BUF_X1 \RegFile/_8499_ ( .A(\RegFile/reg_0 [6] ), .Z(\RegFile/_3310_ ) );
BUF_X1 \RegFile/_8500_ ( .A(\RegFile/_0058_ ), .Z(\RegFile/_0122_ ) );
BUF_X1 \RegFile/_8501_ ( .A(\RegFile/_0676_ ), .Z(\_RegFile_io_rd1 [6] ) );
BUF_X1 \RegFile/_8502_ ( .A(\RegFile/_0061_ ), .Z(\RegFile/_0125_ ) );
BUF_X1 \RegFile/_8503_ ( .A(\RegFile/reg_13 [7] ), .Z(\RegFile/_3439_ ) );
BUF_X1 \RegFile/_8504_ ( .A(\RegFile/reg_12 [7] ), .Z(\RegFile/_3407_ ) );
BUF_X1 \RegFile/_8505_ ( .A(\RegFile/reg_11 [7] ), .Z(\RegFile/_3375_ ) );
BUF_X1 \RegFile/_8506_ ( .A(\RegFile/reg_10 [7] ), .Z(\RegFile/_3343_ ) );
BUF_X1 \RegFile/_8507_ ( .A(\RegFile/reg_9 [7] ), .Z(\RegFile/_3791_ ) );
BUF_X1 \RegFile/_8508_ ( .A(\RegFile/reg_8 [7] ), .Z(\RegFile/_3759_ ) );
BUF_X1 \RegFile/_8509_ ( .A(\RegFile/reg_7 [7] ), .Z(\RegFile/_3727_ ) );
BUF_X1 \RegFile/_8510_ ( .A(\RegFile/reg_6 [7] ), .Z(\RegFile/_3695_ ) );
BUF_X1 \RegFile/_8511_ ( .A(\RegFile/reg_5 [7] ), .Z(\RegFile/_3663_ ) );
BUF_X1 \RegFile/_8512_ ( .A(\RegFile/reg_4 [7] ), .Z(\RegFile/_3631_ ) );
BUF_X1 \RegFile/_8513_ ( .A(\RegFile/reg_3 [7] ), .Z(\RegFile/_3599_ ) );
BUF_X1 \RegFile/_8514_ ( .A(\RegFile/reg_2 [7] ), .Z(\RegFile/_3567_ ) );
BUF_X1 \RegFile/_8515_ ( .A(\RegFile/reg_1 [7] ), .Z(\RegFile/_3535_ ) );
BUF_X1 \RegFile/_8516_ ( .A(\RegFile/reg_0 [7] ), .Z(\RegFile/_3311_ ) );
BUF_X1 \RegFile/_8517_ ( .A(\RegFile/_0060_ ), .Z(\RegFile/_0124_ ) );
BUF_X1 \RegFile/_8518_ ( .A(\RegFile/_0677_ ), .Z(\_RegFile_io_rd1 [7] ) );
BUF_X1 \RegFile/_8519_ ( .A(\RegFile/_0063_ ), .Z(\RegFile/_0127_ ) );
BUF_X1 \RegFile/_8520_ ( .A(\RegFile/reg_13 [8] ), .Z(\RegFile/_3440_ ) );
BUF_X1 \RegFile/_8521_ ( .A(\RegFile/reg_12 [8] ), .Z(\RegFile/_3408_ ) );
BUF_X1 \RegFile/_8522_ ( .A(\RegFile/reg_11 [8] ), .Z(\RegFile/_3376_ ) );
BUF_X1 \RegFile/_8523_ ( .A(\RegFile/reg_10 [8] ), .Z(\RegFile/_3344_ ) );
BUF_X1 \RegFile/_8524_ ( .A(\RegFile/reg_9 [8] ), .Z(\RegFile/_3792_ ) );
BUF_X1 \RegFile/_8525_ ( .A(\RegFile/reg_8 [8] ), .Z(\RegFile/_3760_ ) );
BUF_X1 \RegFile/_8526_ ( .A(\RegFile/reg_7 [8] ), .Z(\RegFile/_3728_ ) );
BUF_X1 \RegFile/_8527_ ( .A(\RegFile/reg_6 [8] ), .Z(\RegFile/_3696_ ) );
BUF_X1 \RegFile/_8528_ ( .A(\RegFile/reg_5 [8] ), .Z(\RegFile/_3664_ ) );
BUF_X1 \RegFile/_8529_ ( .A(\RegFile/reg_4 [8] ), .Z(\RegFile/_3632_ ) );
BUF_X1 \RegFile/_8530_ ( .A(\RegFile/reg_3 [8] ), .Z(\RegFile/_3600_ ) );
BUF_X1 \RegFile/_8531_ ( .A(\RegFile/reg_2 [8] ), .Z(\RegFile/_3568_ ) );
BUF_X1 \RegFile/_8532_ ( .A(\RegFile/reg_1 [8] ), .Z(\RegFile/_3536_ ) );
BUF_X1 \RegFile/_8533_ ( .A(\RegFile/reg_0 [8] ), .Z(\RegFile/_3312_ ) );
BUF_X1 \RegFile/_8534_ ( .A(\RegFile/_0062_ ), .Z(\RegFile/_0126_ ) );
BUF_X1 \RegFile/_8535_ ( .A(\RegFile/_0678_ ), .Z(\_RegFile_io_rd1 [8] ) );
BUF_X1 \RegFile/_8536_ ( .A(\RegFile/_0001_ ), .Z(\RegFile/_0065_ ) );
BUF_X1 \RegFile/_8537_ ( .A(\RegFile/reg_13 [9] ), .Z(\RegFile/_3441_ ) );
BUF_X1 \RegFile/_8538_ ( .A(\RegFile/reg_12 [9] ), .Z(\RegFile/_3409_ ) );
BUF_X1 \RegFile/_8539_ ( .A(\RegFile/reg_11 [9] ), .Z(\RegFile/_3377_ ) );
BUF_X1 \RegFile/_8540_ ( .A(\RegFile/reg_10 [9] ), .Z(\RegFile/_3345_ ) );
BUF_X1 \RegFile/_8541_ ( .A(\RegFile/reg_9 [9] ), .Z(\RegFile/_3793_ ) );
BUF_X1 \RegFile/_8542_ ( .A(\RegFile/reg_8 [9] ), .Z(\RegFile/_3761_ ) );
BUF_X1 \RegFile/_8543_ ( .A(\RegFile/reg_7 [9] ), .Z(\RegFile/_3729_ ) );
BUF_X1 \RegFile/_8544_ ( .A(\RegFile/reg_6 [9] ), .Z(\RegFile/_3697_ ) );
BUF_X1 \RegFile/_8545_ ( .A(\RegFile/reg_5 [9] ), .Z(\RegFile/_3665_ ) );
BUF_X1 \RegFile/_8546_ ( .A(\RegFile/reg_4 [9] ), .Z(\RegFile/_3633_ ) );
BUF_X1 \RegFile/_8547_ ( .A(\RegFile/reg_3 [9] ), .Z(\RegFile/_3601_ ) );
BUF_X1 \RegFile/_8548_ ( .A(\RegFile/reg_2 [9] ), .Z(\RegFile/_3569_ ) );
BUF_X1 \RegFile/_8549_ ( .A(\RegFile/reg_1 [9] ), .Z(\RegFile/_3537_ ) );
BUF_X1 \RegFile/_8550_ ( .A(\RegFile/reg_0 [9] ), .Z(\RegFile/_3313_ ) );
BUF_X1 \RegFile/_8551_ ( .A(\RegFile/_0000_ ), .Z(\RegFile/_0064_ ) );
BUF_X1 \RegFile/_8552_ ( .A(\RegFile/_0679_ ), .Z(\_RegFile_io_rd1 [9] ) );
BUF_X1 \RegFile/_8553_ ( .A(\RegFile/_0003_ ), .Z(\RegFile/_0067_ ) );
BUF_X1 \RegFile/_8554_ ( .A(\RegFile/reg_13 [10] ), .Z(\RegFile/_3411_ ) );
BUF_X1 \RegFile/_8555_ ( .A(\RegFile/reg_12 [10] ), .Z(\RegFile/_3379_ ) );
BUF_X1 \RegFile/_8556_ ( .A(\RegFile/reg_11 [10] ), .Z(\RegFile/_3347_ ) );
BUF_X1 \RegFile/_8557_ ( .A(\RegFile/reg_10 [10] ), .Z(\RegFile/_3315_ ) );
BUF_X1 \RegFile/_8558_ ( .A(\RegFile/reg_9 [10] ), .Z(\RegFile/_3763_ ) );
BUF_X1 \RegFile/_8559_ ( .A(\RegFile/reg_8 [10] ), .Z(\RegFile/_3731_ ) );
BUF_X1 \RegFile/_8560_ ( .A(\RegFile/reg_7 [10] ), .Z(\RegFile/_3699_ ) );
BUF_X1 \RegFile/_8561_ ( .A(\RegFile/reg_6 [10] ), .Z(\RegFile/_3667_ ) );
BUF_X1 \RegFile/_8562_ ( .A(\RegFile/reg_5 [10] ), .Z(\RegFile/_3635_ ) );
BUF_X1 \RegFile/_8563_ ( .A(\RegFile/reg_4 [10] ), .Z(\RegFile/_3603_ ) );
BUF_X1 \RegFile/_8564_ ( .A(\RegFile/reg_3 [10] ), .Z(\RegFile/_3571_ ) );
BUF_X1 \RegFile/_8565_ ( .A(\RegFile/reg_2 [10] ), .Z(\RegFile/_3539_ ) );
BUF_X1 \RegFile/_8566_ ( .A(\RegFile/reg_1 [10] ), .Z(\RegFile/_3507_ ) );
BUF_X1 \RegFile/_8567_ ( .A(\RegFile/reg_0 [10] ), .Z(\RegFile/_3283_ ) );
BUF_X1 \RegFile/_8568_ ( .A(\RegFile/_0002_ ), .Z(\RegFile/_0066_ ) );
BUF_X1 \RegFile/_8569_ ( .A(\RegFile/_0649_ ), .Z(\_RegFile_io_rd1 [10] ) );
BUF_X1 \RegFile/_8570_ ( .A(\RegFile/_0005_ ), .Z(\RegFile/_0069_ ) );
BUF_X1 \RegFile/_8571_ ( .A(\RegFile/reg_13 [11] ), .Z(\RegFile/_3412_ ) );
BUF_X1 \RegFile/_8572_ ( .A(\RegFile/reg_12 [11] ), .Z(\RegFile/_3380_ ) );
BUF_X1 \RegFile/_8573_ ( .A(\RegFile/reg_11 [11] ), .Z(\RegFile/_3348_ ) );
BUF_X1 \RegFile/_8574_ ( .A(\RegFile/reg_10 [11] ), .Z(\RegFile/_3316_ ) );
BUF_X1 \RegFile/_8575_ ( .A(\RegFile/reg_9 [11] ), .Z(\RegFile/_3764_ ) );
BUF_X1 \RegFile/_8576_ ( .A(\RegFile/reg_8 [11] ), .Z(\RegFile/_3732_ ) );
BUF_X1 \RegFile/_8577_ ( .A(\RegFile/reg_7 [11] ), .Z(\RegFile/_3700_ ) );
BUF_X1 \RegFile/_8578_ ( .A(\RegFile/reg_6 [11] ), .Z(\RegFile/_3668_ ) );
BUF_X1 \RegFile/_8579_ ( .A(\RegFile/reg_5 [11] ), .Z(\RegFile/_3636_ ) );
BUF_X1 \RegFile/_8580_ ( .A(\RegFile/reg_4 [11] ), .Z(\RegFile/_3604_ ) );
BUF_X1 \RegFile/_8581_ ( .A(\RegFile/reg_3 [11] ), .Z(\RegFile/_3572_ ) );
BUF_X1 \RegFile/_8582_ ( .A(\RegFile/reg_2 [11] ), .Z(\RegFile/_3540_ ) );
BUF_X1 \RegFile/_8583_ ( .A(\RegFile/reg_1 [11] ), .Z(\RegFile/_3508_ ) );
BUF_X1 \RegFile/_8584_ ( .A(\RegFile/reg_0 [11] ), .Z(\RegFile/_3284_ ) );
BUF_X1 \RegFile/_8585_ ( .A(\RegFile/_0004_ ), .Z(\RegFile/_0068_ ) );
BUF_X1 \RegFile/_8586_ ( .A(\RegFile/_0650_ ), .Z(\_RegFile_io_rd1 [11] ) );
BUF_X1 \RegFile/_8587_ ( .A(\RegFile/_0007_ ), .Z(\RegFile/_0071_ ) );
BUF_X1 \RegFile/_8588_ ( .A(\RegFile/reg_13 [12] ), .Z(\RegFile/_3413_ ) );
BUF_X1 \RegFile/_8589_ ( .A(\RegFile/reg_12 [12] ), .Z(\RegFile/_3381_ ) );
BUF_X1 \RegFile/_8590_ ( .A(\RegFile/reg_11 [12] ), .Z(\RegFile/_3349_ ) );
BUF_X1 \RegFile/_8591_ ( .A(\RegFile/reg_10 [12] ), .Z(\RegFile/_3317_ ) );
BUF_X1 \RegFile/_8592_ ( .A(\RegFile/reg_9 [12] ), .Z(\RegFile/_3765_ ) );
BUF_X1 \RegFile/_8593_ ( .A(\RegFile/reg_8 [12] ), .Z(\RegFile/_3733_ ) );
BUF_X1 \RegFile/_8594_ ( .A(\RegFile/reg_7 [12] ), .Z(\RegFile/_3701_ ) );
BUF_X1 \RegFile/_8595_ ( .A(\RegFile/reg_6 [12] ), .Z(\RegFile/_3669_ ) );
BUF_X1 \RegFile/_8596_ ( .A(\RegFile/reg_5 [12] ), .Z(\RegFile/_3637_ ) );
BUF_X1 \RegFile/_8597_ ( .A(\RegFile/reg_4 [12] ), .Z(\RegFile/_3605_ ) );
BUF_X1 \RegFile/_8598_ ( .A(\RegFile/reg_3 [12] ), .Z(\RegFile/_3573_ ) );
BUF_X1 \RegFile/_8599_ ( .A(\RegFile/reg_2 [12] ), .Z(\RegFile/_3541_ ) );
BUF_X1 \RegFile/_8600_ ( .A(\RegFile/reg_1 [12] ), .Z(\RegFile/_3509_ ) );
BUF_X1 \RegFile/_8601_ ( .A(\RegFile/reg_0 [12] ), .Z(\RegFile/_3285_ ) );
BUF_X1 \RegFile/_8602_ ( .A(\RegFile/_0006_ ), .Z(\RegFile/_0070_ ) );
BUF_X1 \RegFile/_8603_ ( .A(\RegFile/_0651_ ), .Z(\_RegFile_io_rd1 [12] ) );
BUF_X1 \RegFile/_8604_ ( .A(\RegFile/_0009_ ), .Z(\RegFile/_0073_ ) );
BUF_X1 \RegFile/_8605_ ( .A(\RegFile/reg_13 [13] ), .Z(\RegFile/_3414_ ) );
BUF_X1 \RegFile/_8606_ ( .A(\RegFile/reg_12 [13] ), .Z(\RegFile/_3382_ ) );
BUF_X1 \RegFile/_8607_ ( .A(\RegFile/reg_11 [13] ), .Z(\RegFile/_3350_ ) );
BUF_X1 \RegFile/_8608_ ( .A(\RegFile/reg_10 [13] ), .Z(\RegFile/_3318_ ) );
BUF_X1 \RegFile/_8609_ ( .A(\RegFile/reg_9 [13] ), .Z(\RegFile/_3766_ ) );
BUF_X1 \RegFile/_8610_ ( .A(\RegFile/reg_8 [13] ), .Z(\RegFile/_3734_ ) );
BUF_X1 \RegFile/_8611_ ( .A(\RegFile/reg_7 [13] ), .Z(\RegFile/_3702_ ) );
BUF_X1 \RegFile/_8612_ ( .A(\RegFile/reg_6 [13] ), .Z(\RegFile/_3670_ ) );
BUF_X1 \RegFile/_8613_ ( .A(\RegFile/reg_5 [13] ), .Z(\RegFile/_3638_ ) );
BUF_X1 \RegFile/_8614_ ( .A(\RegFile/reg_4 [13] ), .Z(\RegFile/_3606_ ) );
BUF_X1 \RegFile/_8615_ ( .A(\RegFile/reg_3 [13] ), .Z(\RegFile/_3574_ ) );
BUF_X1 \RegFile/_8616_ ( .A(\RegFile/reg_2 [13] ), .Z(\RegFile/_3542_ ) );
BUF_X1 \RegFile/_8617_ ( .A(\RegFile/reg_1 [13] ), .Z(\RegFile/_3510_ ) );
BUF_X1 \RegFile/_8618_ ( .A(\RegFile/reg_0 [13] ), .Z(\RegFile/_3286_ ) );
BUF_X1 \RegFile/_8619_ ( .A(\RegFile/_0008_ ), .Z(\RegFile/_0072_ ) );
BUF_X1 \RegFile/_8620_ ( .A(\RegFile/_0652_ ), .Z(\_RegFile_io_rd1 [13] ) );
BUF_X1 \RegFile/_8621_ ( .A(\RegFile/_0011_ ), .Z(\RegFile/_0075_ ) );
BUF_X1 \RegFile/_8622_ ( .A(\RegFile/reg_13 [14] ), .Z(\RegFile/_3415_ ) );
BUF_X1 \RegFile/_8623_ ( .A(\RegFile/reg_12 [14] ), .Z(\RegFile/_3383_ ) );
BUF_X1 \RegFile/_8624_ ( .A(\RegFile/reg_11 [14] ), .Z(\RegFile/_3351_ ) );
BUF_X1 \RegFile/_8625_ ( .A(\RegFile/reg_10 [14] ), .Z(\RegFile/_3319_ ) );
BUF_X1 \RegFile/_8626_ ( .A(\RegFile/reg_9 [14] ), .Z(\RegFile/_3767_ ) );
BUF_X1 \RegFile/_8627_ ( .A(\RegFile/reg_8 [14] ), .Z(\RegFile/_3735_ ) );
BUF_X1 \RegFile/_8628_ ( .A(\RegFile/reg_7 [14] ), .Z(\RegFile/_3703_ ) );
BUF_X1 \RegFile/_8629_ ( .A(\RegFile/reg_6 [14] ), .Z(\RegFile/_3671_ ) );
BUF_X1 \RegFile/_8630_ ( .A(\RegFile/reg_5 [14] ), .Z(\RegFile/_3639_ ) );
BUF_X1 \RegFile/_8631_ ( .A(\RegFile/reg_4 [14] ), .Z(\RegFile/_3607_ ) );
BUF_X1 \RegFile/_8632_ ( .A(\RegFile/reg_3 [14] ), .Z(\RegFile/_3575_ ) );
BUF_X1 \RegFile/_8633_ ( .A(\RegFile/reg_2 [14] ), .Z(\RegFile/_3543_ ) );
BUF_X1 \RegFile/_8634_ ( .A(\RegFile/reg_1 [14] ), .Z(\RegFile/_3511_ ) );
BUF_X1 \RegFile/_8635_ ( .A(\RegFile/reg_0 [14] ), .Z(\RegFile/_3287_ ) );
BUF_X1 \RegFile/_8636_ ( .A(\RegFile/_0010_ ), .Z(\RegFile/_0074_ ) );
BUF_X1 \RegFile/_8637_ ( .A(\RegFile/_0653_ ), .Z(\_RegFile_io_rd1 [14] ) );
BUF_X1 \RegFile/_8638_ ( .A(\RegFile/_0013_ ), .Z(\RegFile/_0077_ ) );
BUF_X1 \RegFile/_8639_ ( .A(\RegFile/reg_13 [15] ), .Z(\RegFile/_3416_ ) );
BUF_X1 \RegFile/_8640_ ( .A(\RegFile/reg_12 [15] ), .Z(\RegFile/_3384_ ) );
BUF_X1 \RegFile/_8641_ ( .A(\RegFile/reg_11 [15] ), .Z(\RegFile/_3352_ ) );
BUF_X1 \RegFile/_8642_ ( .A(\RegFile/reg_10 [15] ), .Z(\RegFile/_3320_ ) );
BUF_X1 \RegFile/_8643_ ( .A(\RegFile/reg_9 [15] ), .Z(\RegFile/_3768_ ) );
BUF_X1 \RegFile/_8644_ ( .A(\RegFile/reg_8 [15] ), .Z(\RegFile/_3736_ ) );
BUF_X1 \RegFile/_8645_ ( .A(\RegFile/reg_7 [15] ), .Z(\RegFile/_3704_ ) );
BUF_X1 \RegFile/_8646_ ( .A(\RegFile/reg_6 [15] ), .Z(\RegFile/_3672_ ) );
BUF_X1 \RegFile/_8647_ ( .A(\RegFile/reg_5 [15] ), .Z(\RegFile/_3640_ ) );
BUF_X1 \RegFile/_8648_ ( .A(\RegFile/reg_4 [15] ), .Z(\RegFile/_3608_ ) );
BUF_X1 \RegFile/_8649_ ( .A(\RegFile/reg_3 [15] ), .Z(\RegFile/_3576_ ) );
BUF_X1 \RegFile/_8650_ ( .A(\RegFile/reg_2 [15] ), .Z(\RegFile/_3544_ ) );
BUF_X1 \RegFile/_8651_ ( .A(\RegFile/reg_1 [15] ), .Z(\RegFile/_3512_ ) );
BUF_X1 \RegFile/_8652_ ( .A(\RegFile/reg_0 [15] ), .Z(\RegFile/_3288_ ) );
BUF_X1 \RegFile/_8653_ ( .A(\RegFile/_0012_ ), .Z(\RegFile/_0076_ ) );
BUF_X1 \RegFile/_8654_ ( .A(\RegFile/_0654_ ), .Z(\_RegFile_io_rd1 [15] ) );
BUF_X1 \RegFile/_8655_ ( .A(\RegFile/_0015_ ), .Z(\RegFile/_0079_ ) );
BUF_X1 \RegFile/_8656_ ( .A(\RegFile/reg_13 [16] ), .Z(\RegFile/_3417_ ) );
BUF_X1 \RegFile/_8657_ ( .A(\RegFile/reg_12 [16] ), .Z(\RegFile/_3385_ ) );
BUF_X1 \RegFile/_8658_ ( .A(\RegFile/reg_11 [16] ), .Z(\RegFile/_3353_ ) );
BUF_X1 \RegFile/_8659_ ( .A(\RegFile/reg_10 [16] ), .Z(\RegFile/_3321_ ) );
BUF_X1 \RegFile/_8660_ ( .A(\RegFile/reg_9 [16] ), .Z(\RegFile/_3769_ ) );
BUF_X1 \RegFile/_8661_ ( .A(\RegFile/reg_8 [16] ), .Z(\RegFile/_3737_ ) );
BUF_X1 \RegFile/_8662_ ( .A(\RegFile/reg_7 [16] ), .Z(\RegFile/_3705_ ) );
BUF_X1 \RegFile/_8663_ ( .A(\RegFile/reg_6 [16] ), .Z(\RegFile/_3673_ ) );
BUF_X1 \RegFile/_8664_ ( .A(\RegFile/reg_5 [16] ), .Z(\RegFile/_3641_ ) );
BUF_X1 \RegFile/_8665_ ( .A(\RegFile/reg_4 [16] ), .Z(\RegFile/_3609_ ) );
BUF_X1 \RegFile/_8666_ ( .A(\RegFile/reg_3 [16] ), .Z(\RegFile/_3577_ ) );
BUF_X1 \RegFile/_8667_ ( .A(\RegFile/reg_2 [16] ), .Z(\RegFile/_3545_ ) );
BUF_X1 \RegFile/_8668_ ( .A(\RegFile/reg_1 [16] ), .Z(\RegFile/_3513_ ) );
BUF_X1 \RegFile/_8669_ ( .A(\RegFile/reg_0 [16] ), .Z(\RegFile/_3289_ ) );
BUF_X1 \RegFile/_8670_ ( .A(\RegFile/_0014_ ), .Z(\RegFile/_0078_ ) );
BUF_X1 \RegFile/_8671_ ( .A(\RegFile/_0655_ ), .Z(\_RegFile_io_rd1 [16] ) );
BUF_X1 \RegFile/_8672_ ( .A(\RegFile/_0017_ ), .Z(\RegFile/_0081_ ) );
BUF_X1 \RegFile/_8673_ ( .A(\RegFile/reg_13 [17] ), .Z(\RegFile/_3418_ ) );
BUF_X1 \RegFile/_8674_ ( .A(\RegFile/reg_12 [17] ), .Z(\RegFile/_3386_ ) );
BUF_X1 \RegFile/_8675_ ( .A(\RegFile/reg_11 [17] ), .Z(\RegFile/_3354_ ) );
BUF_X1 \RegFile/_8676_ ( .A(\RegFile/reg_10 [17] ), .Z(\RegFile/_3322_ ) );
BUF_X1 \RegFile/_8677_ ( .A(\RegFile/reg_9 [17] ), .Z(\RegFile/_3770_ ) );
BUF_X1 \RegFile/_8678_ ( .A(\RegFile/reg_8 [17] ), .Z(\RegFile/_3738_ ) );
BUF_X1 \RegFile/_8679_ ( .A(\RegFile/reg_7 [17] ), .Z(\RegFile/_3706_ ) );
BUF_X1 \RegFile/_8680_ ( .A(\RegFile/reg_6 [17] ), .Z(\RegFile/_3674_ ) );
BUF_X1 \RegFile/_8681_ ( .A(\RegFile/reg_5 [17] ), .Z(\RegFile/_3642_ ) );
BUF_X1 \RegFile/_8682_ ( .A(\RegFile/reg_4 [17] ), .Z(\RegFile/_3610_ ) );
BUF_X1 \RegFile/_8683_ ( .A(\RegFile/reg_3 [17] ), .Z(\RegFile/_3578_ ) );
BUF_X1 \RegFile/_8684_ ( .A(\RegFile/reg_2 [17] ), .Z(\RegFile/_3546_ ) );
BUF_X1 \RegFile/_8685_ ( .A(\RegFile/reg_1 [17] ), .Z(\RegFile/_3514_ ) );
BUF_X1 \RegFile/_8686_ ( .A(\RegFile/reg_0 [17] ), .Z(\RegFile/_3290_ ) );
BUF_X1 \RegFile/_8687_ ( .A(\RegFile/_0016_ ), .Z(\RegFile/_0080_ ) );
BUF_X1 \RegFile/_8688_ ( .A(\RegFile/_0656_ ), .Z(\_RegFile_io_rd1 [17] ) );
BUF_X1 \RegFile/_8689_ ( .A(\RegFile/_0019_ ), .Z(\RegFile/_0083_ ) );
BUF_X1 \RegFile/_8690_ ( .A(\RegFile/reg_13 [18] ), .Z(\RegFile/_3419_ ) );
BUF_X1 \RegFile/_8691_ ( .A(\RegFile/reg_12 [18] ), .Z(\RegFile/_3387_ ) );
BUF_X1 \RegFile/_8692_ ( .A(\RegFile/reg_11 [18] ), .Z(\RegFile/_3355_ ) );
BUF_X1 \RegFile/_8693_ ( .A(\RegFile/reg_10 [18] ), .Z(\RegFile/_3323_ ) );
BUF_X1 \RegFile/_8694_ ( .A(\RegFile/reg_9 [18] ), .Z(\RegFile/_3771_ ) );
BUF_X1 \RegFile/_8695_ ( .A(\RegFile/reg_8 [18] ), .Z(\RegFile/_3739_ ) );
BUF_X1 \RegFile/_8696_ ( .A(\RegFile/reg_7 [18] ), .Z(\RegFile/_3707_ ) );
BUF_X1 \RegFile/_8697_ ( .A(\RegFile/reg_6 [18] ), .Z(\RegFile/_3675_ ) );
BUF_X1 \RegFile/_8698_ ( .A(\RegFile/reg_5 [18] ), .Z(\RegFile/_3643_ ) );
BUF_X1 \RegFile/_8699_ ( .A(\RegFile/reg_4 [18] ), .Z(\RegFile/_3611_ ) );
BUF_X1 \RegFile/_8700_ ( .A(\RegFile/reg_3 [18] ), .Z(\RegFile/_3579_ ) );
BUF_X1 \RegFile/_8701_ ( .A(\RegFile/reg_2 [18] ), .Z(\RegFile/_3547_ ) );
BUF_X1 \RegFile/_8702_ ( .A(\RegFile/reg_1 [18] ), .Z(\RegFile/_3515_ ) );
BUF_X1 \RegFile/_8703_ ( .A(\RegFile/reg_0 [18] ), .Z(\RegFile/_3291_ ) );
BUF_X1 \RegFile/_8704_ ( .A(\RegFile/_0018_ ), .Z(\RegFile/_0082_ ) );
BUF_X1 \RegFile/_8705_ ( .A(\RegFile/_0657_ ), .Z(\_RegFile_io_rd1 [18] ) );
BUF_X1 \RegFile/_8706_ ( .A(\RegFile/_0021_ ), .Z(\RegFile/_0085_ ) );
BUF_X1 \RegFile/_8707_ ( .A(\RegFile/reg_13 [19] ), .Z(\RegFile/_3420_ ) );
BUF_X1 \RegFile/_8708_ ( .A(\RegFile/reg_12 [19] ), .Z(\RegFile/_3388_ ) );
BUF_X1 \RegFile/_8709_ ( .A(\RegFile/reg_11 [19] ), .Z(\RegFile/_3356_ ) );
BUF_X1 \RegFile/_8710_ ( .A(\RegFile/reg_10 [19] ), .Z(\RegFile/_3324_ ) );
BUF_X1 \RegFile/_8711_ ( .A(\RegFile/reg_9 [19] ), .Z(\RegFile/_3772_ ) );
BUF_X1 \RegFile/_8712_ ( .A(\RegFile/reg_8 [19] ), .Z(\RegFile/_3740_ ) );
BUF_X1 \RegFile/_8713_ ( .A(\RegFile/reg_7 [19] ), .Z(\RegFile/_3708_ ) );
BUF_X1 \RegFile/_8714_ ( .A(\RegFile/reg_6 [19] ), .Z(\RegFile/_3676_ ) );
BUF_X1 \RegFile/_8715_ ( .A(\RegFile/reg_5 [19] ), .Z(\RegFile/_3644_ ) );
BUF_X1 \RegFile/_8716_ ( .A(\RegFile/reg_4 [19] ), .Z(\RegFile/_3612_ ) );
BUF_X1 \RegFile/_8717_ ( .A(\RegFile/reg_3 [19] ), .Z(\RegFile/_3580_ ) );
BUF_X1 \RegFile/_8718_ ( .A(\RegFile/reg_2 [19] ), .Z(\RegFile/_3548_ ) );
BUF_X1 \RegFile/_8719_ ( .A(\RegFile/reg_1 [19] ), .Z(\RegFile/_3516_ ) );
BUF_X1 \RegFile/_8720_ ( .A(\RegFile/reg_0 [19] ), .Z(\RegFile/_3292_ ) );
BUF_X1 \RegFile/_8721_ ( .A(\RegFile/_0020_ ), .Z(\RegFile/_0084_ ) );
BUF_X1 \RegFile/_8722_ ( .A(\RegFile/_0658_ ), .Z(\_RegFile_io_rd1 [19] ) );
BUF_X1 \RegFile/_8723_ ( .A(\RegFile/_0023_ ), .Z(\RegFile/_0087_ ) );
BUF_X1 \RegFile/_8724_ ( .A(\RegFile/reg_13 [20] ), .Z(\RegFile/_3422_ ) );
BUF_X1 \RegFile/_8725_ ( .A(\RegFile/reg_12 [20] ), .Z(\RegFile/_3390_ ) );
BUF_X1 \RegFile/_8726_ ( .A(\RegFile/reg_11 [20] ), .Z(\RegFile/_3358_ ) );
BUF_X1 \RegFile/_8727_ ( .A(\RegFile/reg_10 [20] ), .Z(\RegFile/_3326_ ) );
BUF_X1 \RegFile/_8728_ ( .A(\RegFile/reg_9 [20] ), .Z(\RegFile/_3774_ ) );
BUF_X1 \RegFile/_8729_ ( .A(\RegFile/reg_8 [20] ), .Z(\RegFile/_3742_ ) );
BUF_X1 \RegFile/_8730_ ( .A(\RegFile/reg_7 [20] ), .Z(\RegFile/_3710_ ) );
BUF_X1 \RegFile/_8731_ ( .A(\RegFile/reg_6 [20] ), .Z(\RegFile/_3678_ ) );
BUF_X1 \RegFile/_8732_ ( .A(\RegFile/reg_5 [20] ), .Z(\RegFile/_3646_ ) );
BUF_X1 \RegFile/_8733_ ( .A(\RegFile/reg_4 [20] ), .Z(\RegFile/_3614_ ) );
BUF_X1 \RegFile/_8734_ ( .A(\RegFile/reg_3 [20] ), .Z(\RegFile/_3582_ ) );
BUF_X1 \RegFile/_8735_ ( .A(\RegFile/reg_2 [20] ), .Z(\RegFile/_3550_ ) );
BUF_X1 \RegFile/_8736_ ( .A(\RegFile/reg_1 [20] ), .Z(\RegFile/_3518_ ) );
BUF_X1 \RegFile/_8737_ ( .A(\RegFile/reg_0 [20] ), .Z(\RegFile/_3294_ ) );
BUF_X1 \RegFile/_8738_ ( .A(\RegFile/_0022_ ), .Z(\RegFile/_0086_ ) );
BUF_X1 \RegFile/_8739_ ( .A(\RegFile/_0660_ ), .Z(\_RegFile_io_rd1 [20] ) );
BUF_X1 \RegFile/_8740_ ( .A(\RegFile/_0025_ ), .Z(\RegFile/_0089_ ) );
BUF_X1 \RegFile/_8741_ ( .A(\RegFile/reg_13 [21] ), .Z(\RegFile/_3423_ ) );
BUF_X1 \RegFile/_8742_ ( .A(\RegFile/reg_12 [21] ), .Z(\RegFile/_3391_ ) );
BUF_X1 \RegFile/_8743_ ( .A(\RegFile/reg_11 [21] ), .Z(\RegFile/_3359_ ) );
BUF_X1 \RegFile/_8744_ ( .A(\RegFile/reg_10 [21] ), .Z(\RegFile/_3327_ ) );
BUF_X1 \RegFile/_8745_ ( .A(\RegFile/reg_9 [21] ), .Z(\RegFile/_3775_ ) );
BUF_X1 \RegFile/_8746_ ( .A(\RegFile/reg_8 [21] ), .Z(\RegFile/_3743_ ) );
BUF_X1 \RegFile/_8747_ ( .A(\RegFile/reg_7 [21] ), .Z(\RegFile/_3711_ ) );
BUF_X1 \RegFile/_8748_ ( .A(\RegFile/reg_6 [21] ), .Z(\RegFile/_3679_ ) );
BUF_X1 \RegFile/_8749_ ( .A(\RegFile/reg_5 [21] ), .Z(\RegFile/_3647_ ) );
BUF_X1 \RegFile/_8750_ ( .A(\RegFile/reg_4 [21] ), .Z(\RegFile/_3615_ ) );
BUF_X1 \RegFile/_8751_ ( .A(\RegFile/reg_3 [21] ), .Z(\RegFile/_3583_ ) );
BUF_X1 \RegFile/_8752_ ( .A(\RegFile/reg_2 [21] ), .Z(\RegFile/_3551_ ) );
BUF_X1 \RegFile/_8753_ ( .A(\RegFile/reg_1 [21] ), .Z(\RegFile/_3519_ ) );
BUF_X1 \RegFile/_8754_ ( .A(\RegFile/reg_0 [21] ), .Z(\RegFile/_3295_ ) );
BUF_X1 \RegFile/_8755_ ( .A(\RegFile/_0024_ ), .Z(\RegFile/_0088_ ) );
BUF_X1 \RegFile/_8756_ ( .A(\RegFile/_0661_ ), .Z(\_RegFile_io_rd1 [21] ) );
BUF_X1 \RegFile/_8757_ ( .A(\RegFile/_0027_ ), .Z(\RegFile/_0091_ ) );
BUF_X1 \RegFile/_8758_ ( .A(\RegFile/reg_13 [22] ), .Z(\RegFile/_3424_ ) );
BUF_X1 \RegFile/_8759_ ( .A(\RegFile/reg_12 [22] ), .Z(\RegFile/_3392_ ) );
BUF_X1 \RegFile/_8760_ ( .A(\RegFile/reg_11 [22] ), .Z(\RegFile/_3360_ ) );
BUF_X1 \RegFile/_8761_ ( .A(\RegFile/reg_10 [22] ), .Z(\RegFile/_3328_ ) );
BUF_X1 \RegFile/_8762_ ( .A(\RegFile/reg_9 [22] ), .Z(\RegFile/_3776_ ) );
BUF_X1 \RegFile/_8763_ ( .A(\RegFile/reg_8 [22] ), .Z(\RegFile/_3744_ ) );
BUF_X1 \RegFile/_8764_ ( .A(\RegFile/reg_7 [22] ), .Z(\RegFile/_3712_ ) );
BUF_X1 \RegFile/_8765_ ( .A(\RegFile/reg_6 [22] ), .Z(\RegFile/_3680_ ) );
BUF_X1 \RegFile/_8766_ ( .A(\RegFile/reg_5 [22] ), .Z(\RegFile/_3648_ ) );
BUF_X1 \RegFile/_8767_ ( .A(\RegFile/reg_4 [22] ), .Z(\RegFile/_3616_ ) );
BUF_X1 \RegFile/_8768_ ( .A(\RegFile/reg_3 [22] ), .Z(\RegFile/_3584_ ) );
BUF_X1 \RegFile/_8769_ ( .A(\RegFile/reg_2 [22] ), .Z(\RegFile/_3552_ ) );
BUF_X1 \RegFile/_8770_ ( .A(\RegFile/reg_1 [22] ), .Z(\RegFile/_3520_ ) );
BUF_X1 \RegFile/_8771_ ( .A(\RegFile/reg_0 [22] ), .Z(\RegFile/_3296_ ) );
BUF_X1 \RegFile/_8772_ ( .A(\RegFile/_0026_ ), .Z(\RegFile/_0090_ ) );
BUF_X1 \RegFile/_8773_ ( .A(\RegFile/_0662_ ), .Z(\_RegFile_io_rd1 [22] ) );
BUF_X1 \RegFile/_8774_ ( .A(\RegFile/_0029_ ), .Z(\RegFile/_0093_ ) );
BUF_X1 \RegFile/_8775_ ( .A(\RegFile/reg_13 [23] ), .Z(\RegFile/_3425_ ) );
BUF_X1 \RegFile/_8776_ ( .A(\RegFile/reg_12 [23] ), .Z(\RegFile/_3393_ ) );
BUF_X1 \RegFile/_8777_ ( .A(\RegFile/reg_11 [23] ), .Z(\RegFile/_3361_ ) );
BUF_X1 \RegFile/_8778_ ( .A(\RegFile/reg_10 [23] ), .Z(\RegFile/_3329_ ) );
BUF_X1 \RegFile/_8779_ ( .A(\RegFile/reg_9 [23] ), .Z(\RegFile/_3777_ ) );
BUF_X1 \RegFile/_8780_ ( .A(\RegFile/reg_8 [23] ), .Z(\RegFile/_3745_ ) );
BUF_X1 \RegFile/_8781_ ( .A(\RegFile/reg_7 [23] ), .Z(\RegFile/_3713_ ) );
BUF_X1 \RegFile/_8782_ ( .A(\RegFile/reg_6 [23] ), .Z(\RegFile/_3681_ ) );
BUF_X1 \RegFile/_8783_ ( .A(\RegFile/reg_5 [23] ), .Z(\RegFile/_3649_ ) );
BUF_X1 \RegFile/_8784_ ( .A(\RegFile/reg_4 [23] ), .Z(\RegFile/_3617_ ) );
BUF_X1 \RegFile/_8785_ ( .A(\RegFile/reg_3 [23] ), .Z(\RegFile/_3585_ ) );
BUF_X1 \RegFile/_8786_ ( .A(\RegFile/reg_2 [23] ), .Z(\RegFile/_3553_ ) );
BUF_X1 \RegFile/_8787_ ( .A(\RegFile/reg_1 [23] ), .Z(\RegFile/_3521_ ) );
BUF_X1 \RegFile/_8788_ ( .A(\RegFile/reg_0 [23] ), .Z(\RegFile/_3297_ ) );
BUF_X1 \RegFile/_8789_ ( .A(\RegFile/_0028_ ), .Z(\RegFile/_0092_ ) );
BUF_X1 \RegFile/_8790_ ( .A(\RegFile/_0663_ ), .Z(\_RegFile_io_rd1 [23] ) );
BUF_X1 \RegFile/_8791_ ( .A(\RegFile/_0031_ ), .Z(\RegFile/_0095_ ) );
BUF_X1 \RegFile/_8792_ ( .A(\RegFile/reg_13 [24] ), .Z(\RegFile/_3426_ ) );
BUF_X1 \RegFile/_8793_ ( .A(\RegFile/reg_12 [24] ), .Z(\RegFile/_3394_ ) );
BUF_X1 \RegFile/_8794_ ( .A(\RegFile/reg_11 [24] ), .Z(\RegFile/_3362_ ) );
BUF_X1 \RegFile/_8795_ ( .A(\RegFile/reg_10 [24] ), .Z(\RegFile/_3330_ ) );
BUF_X1 \RegFile/_8796_ ( .A(\RegFile/reg_9 [24] ), .Z(\RegFile/_3778_ ) );
BUF_X1 \RegFile/_8797_ ( .A(\RegFile/reg_8 [24] ), .Z(\RegFile/_3746_ ) );
BUF_X1 \RegFile/_8798_ ( .A(\RegFile/reg_7 [24] ), .Z(\RegFile/_3714_ ) );
BUF_X1 \RegFile/_8799_ ( .A(\RegFile/reg_6 [24] ), .Z(\RegFile/_3682_ ) );
BUF_X1 \RegFile/_8800_ ( .A(\RegFile/reg_5 [24] ), .Z(\RegFile/_3650_ ) );
BUF_X1 \RegFile/_8801_ ( .A(\RegFile/reg_4 [24] ), .Z(\RegFile/_3618_ ) );
BUF_X1 \RegFile/_8802_ ( .A(\RegFile/reg_3 [24] ), .Z(\RegFile/_3586_ ) );
BUF_X1 \RegFile/_8803_ ( .A(\RegFile/reg_2 [24] ), .Z(\RegFile/_3554_ ) );
BUF_X1 \RegFile/_8804_ ( .A(\RegFile/reg_1 [24] ), .Z(\RegFile/_3522_ ) );
BUF_X1 \RegFile/_8805_ ( .A(\RegFile/reg_0 [24] ), .Z(\RegFile/_3298_ ) );
BUF_X1 \RegFile/_8806_ ( .A(\RegFile/_0030_ ), .Z(\RegFile/_0094_ ) );
BUF_X1 \RegFile/_8807_ ( .A(\RegFile/_0664_ ), .Z(\_RegFile_io_rd1 [24] ) );
BUF_X1 \RegFile/_8808_ ( .A(\RegFile/_0033_ ), .Z(\RegFile/_0097_ ) );
BUF_X1 \RegFile/_8809_ ( .A(\RegFile/reg_13 [25] ), .Z(\RegFile/_3427_ ) );
BUF_X1 \RegFile/_8810_ ( .A(\RegFile/reg_12 [25] ), .Z(\RegFile/_3395_ ) );
BUF_X1 \RegFile/_8811_ ( .A(\RegFile/reg_11 [25] ), .Z(\RegFile/_3363_ ) );
BUF_X1 \RegFile/_8812_ ( .A(\RegFile/reg_10 [25] ), .Z(\RegFile/_3331_ ) );
BUF_X1 \RegFile/_8813_ ( .A(\RegFile/reg_9 [25] ), .Z(\RegFile/_3779_ ) );
BUF_X1 \RegFile/_8814_ ( .A(\RegFile/reg_8 [25] ), .Z(\RegFile/_3747_ ) );
BUF_X1 \RegFile/_8815_ ( .A(\RegFile/reg_7 [25] ), .Z(\RegFile/_3715_ ) );
BUF_X1 \RegFile/_8816_ ( .A(\RegFile/reg_6 [25] ), .Z(\RegFile/_3683_ ) );
BUF_X1 \RegFile/_8817_ ( .A(\RegFile/reg_5 [25] ), .Z(\RegFile/_3651_ ) );
BUF_X1 \RegFile/_8818_ ( .A(\RegFile/reg_4 [25] ), .Z(\RegFile/_3619_ ) );
BUF_X1 \RegFile/_8819_ ( .A(\RegFile/reg_3 [25] ), .Z(\RegFile/_3587_ ) );
BUF_X1 \RegFile/_8820_ ( .A(\RegFile/reg_2 [25] ), .Z(\RegFile/_3555_ ) );
BUF_X1 \RegFile/_8821_ ( .A(\RegFile/reg_1 [25] ), .Z(\RegFile/_3523_ ) );
BUF_X1 \RegFile/_8822_ ( .A(\RegFile/reg_0 [25] ), .Z(\RegFile/_3299_ ) );
BUF_X1 \RegFile/_8823_ ( .A(\RegFile/_0032_ ), .Z(\RegFile/_0096_ ) );
BUF_X1 \RegFile/_8824_ ( .A(\RegFile/_0665_ ), .Z(\_RegFile_io_rd1 [25] ) );
BUF_X1 \RegFile/_8825_ ( .A(\RegFile/_0035_ ), .Z(\RegFile/_0099_ ) );
BUF_X1 \RegFile/_8826_ ( .A(\RegFile/reg_13 [26] ), .Z(\RegFile/_3428_ ) );
BUF_X1 \RegFile/_8827_ ( .A(\RegFile/reg_12 [26] ), .Z(\RegFile/_3396_ ) );
BUF_X1 \RegFile/_8828_ ( .A(\RegFile/reg_11 [26] ), .Z(\RegFile/_3364_ ) );
BUF_X1 \RegFile/_8829_ ( .A(\RegFile/reg_10 [26] ), .Z(\RegFile/_3332_ ) );
BUF_X1 \RegFile/_8830_ ( .A(\RegFile/reg_9 [26] ), .Z(\RegFile/_3780_ ) );
BUF_X1 \RegFile/_8831_ ( .A(\RegFile/reg_8 [26] ), .Z(\RegFile/_3748_ ) );
BUF_X1 \RegFile/_8832_ ( .A(\RegFile/reg_7 [26] ), .Z(\RegFile/_3716_ ) );
BUF_X1 \RegFile/_8833_ ( .A(\RegFile/reg_6 [26] ), .Z(\RegFile/_3684_ ) );
BUF_X1 \RegFile/_8834_ ( .A(\RegFile/reg_5 [26] ), .Z(\RegFile/_3652_ ) );
BUF_X1 \RegFile/_8835_ ( .A(\RegFile/reg_4 [26] ), .Z(\RegFile/_3620_ ) );
BUF_X1 \RegFile/_8836_ ( .A(\RegFile/reg_3 [26] ), .Z(\RegFile/_3588_ ) );
BUF_X1 \RegFile/_8837_ ( .A(\RegFile/reg_2 [26] ), .Z(\RegFile/_3556_ ) );
BUF_X1 \RegFile/_8838_ ( .A(\RegFile/reg_1 [26] ), .Z(\RegFile/_3524_ ) );
BUF_X1 \RegFile/_8839_ ( .A(\RegFile/reg_0 [26] ), .Z(\RegFile/_3300_ ) );
BUF_X1 \RegFile/_8840_ ( .A(\RegFile/_0034_ ), .Z(\RegFile/_0098_ ) );
BUF_X1 \RegFile/_8841_ ( .A(\RegFile/_0666_ ), .Z(\_RegFile_io_rd1 [26] ) );
BUF_X1 \RegFile/_8842_ ( .A(\RegFile/_0037_ ), .Z(\RegFile/_0101_ ) );
BUF_X1 \RegFile/_8843_ ( .A(\RegFile/reg_13 [27] ), .Z(\RegFile/_3429_ ) );
BUF_X1 \RegFile/_8844_ ( .A(\RegFile/reg_12 [27] ), .Z(\RegFile/_3397_ ) );
BUF_X1 \RegFile/_8845_ ( .A(\RegFile/reg_11 [27] ), .Z(\RegFile/_3365_ ) );
BUF_X1 \RegFile/_8846_ ( .A(\RegFile/reg_10 [27] ), .Z(\RegFile/_3333_ ) );
BUF_X1 \RegFile/_8847_ ( .A(\RegFile/reg_9 [27] ), .Z(\RegFile/_3781_ ) );
BUF_X1 \RegFile/_8848_ ( .A(\RegFile/reg_8 [27] ), .Z(\RegFile/_3749_ ) );
BUF_X1 \RegFile/_8849_ ( .A(\RegFile/reg_7 [27] ), .Z(\RegFile/_3717_ ) );
BUF_X1 \RegFile/_8850_ ( .A(\RegFile/reg_6 [27] ), .Z(\RegFile/_3685_ ) );
BUF_X1 \RegFile/_8851_ ( .A(\RegFile/reg_5 [27] ), .Z(\RegFile/_3653_ ) );
BUF_X1 \RegFile/_8852_ ( .A(\RegFile/reg_4 [27] ), .Z(\RegFile/_3621_ ) );
BUF_X1 \RegFile/_8853_ ( .A(\RegFile/reg_3 [27] ), .Z(\RegFile/_3589_ ) );
BUF_X1 \RegFile/_8854_ ( .A(\RegFile/reg_2 [27] ), .Z(\RegFile/_3557_ ) );
BUF_X1 \RegFile/_8855_ ( .A(\RegFile/reg_1 [27] ), .Z(\RegFile/_3525_ ) );
BUF_X1 \RegFile/_8856_ ( .A(\RegFile/reg_0 [27] ), .Z(\RegFile/_3301_ ) );
BUF_X1 \RegFile/_8857_ ( .A(\RegFile/_0036_ ), .Z(\RegFile/_0100_ ) );
BUF_X1 \RegFile/_8858_ ( .A(\RegFile/_0667_ ), .Z(\_RegFile_io_rd1 [27] ) );
BUF_X1 \RegFile/_8859_ ( .A(\RegFile/_0039_ ), .Z(\RegFile/_0103_ ) );
BUF_X1 \RegFile/_8860_ ( .A(\RegFile/reg_13 [28] ), .Z(\RegFile/_3430_ ) );
BUF_X1 \RegFile/_8861_ ( .A(\RegFile/reg_12 [28] ), .Z(\RegFile/_3398_ ) );
BUF_X1 \RegFile/_8862_ ( .A(\RegFile/reg_11 [28] ), .Z(\RegFile/_3366_ ) );
BUF_X1 \RegFile/_8863_ ( .A(\RegFile/reg_10 [28] ), .Z(\RegFile/_3334_ ) );
BUF_X1 \RegFile/_8864_ ( .A(\RegFile/reg_9 [28] ), .Z(\RegFile/_3782_ ) );
BUF_X1 \RegFile/_8865_ ( .A(\RegFile/reg_8 [28] ), .Z(\RegFile/_3750_ ) );
BUF_X1 \RegFile/_8866_ ( .A(\RegFile/reg_7 [28] ), .Z(\RegFile/_3718_ ) );
BUF_X1 \RegFile/_8867_ ( .A(\RegFile/reg_6 [28] ), .Z(\RegFile/_3686_ ) );
BUF_X1 \RegFile/_8868_ ( .A(\RegFile/reg_5 [28] ), .Z(\RegFile/_3654_ ) );
BUF_X1 \RegFile/_8869_ ( .A(\RegFile/reg_4 [28] ), .Z(\RegFile/_3622_ ) );
BUF_X1 \RegFile/_8870_ ( .A(\RegFile/reg_3 [28] ), .Z(\RegFile/_3590_ ) );
BUF_X1 \RegFile/_8871_ ( .A(\RegFile/reg_2 [28] ), .Z(\RegFile/_3558_ ) );
BUF_X1 \RegFile/_8872_ ( .A(\RegFile/reg_1 [28] ), .Z(\RegFile/_3526_ ) );
BUF_X1 \RegFile/_8873_ ( .A(\RegFile/reg_0 [28] ), .Z(\RegFile/_3302_ ) );
BUF_X1 \RegFile/_8874_ ( .A(\RegFile/_0038_ ), .Z(\RegFile/_0102_ ) );
BUF_X1 \RegFile/_8875_ ( .A(\RegFile/_0668_ ), .Z(\_RegFile_io_rd1 [28] ) );
BUF_X1 \RegFile/_8876_ ( .A(\RegFile/_0041_ ), .Z(\RegFile/_0105_ ) );
BUF_X1 \RegFile/_8877_ ( .A(\RegFile/reg_13 [29] ), .Z(\RegFile/_3431_ ) );
BUF_X1 \RegFile/_8878_ ( .A(\RegFile/reg_12 [29] ), .Z(\RegFile/_3399_ ) );
BUF_X1 \RegFile/_8879_ ( .A(\RegFile/reg_11 [29] ), .Z(\RegFile/_3367_ ) );
BUF_X1 \RegFile/_8880_ ( .A(\RegFile/reg_10 [29] ), .Z(\RegFile/_3335_ ) );
BUF_X1 \RegFile/_8881_ ( .A(\RegFile/reg_9 [29] ), .Z(\RegFile/_3783_ ) );
BUF_X1 \RegFile/_8882_ ( .A(\RegFile/reg_8 [29] ), .Z(\RegFile/_3751_ ) );
BUF_X1 \RegFile/_8883_ ( .A(\RegFile/reg_7 [29] ), .Z(\RegFile/_3719_ ) );
BUF_X1 \RegFile/_8884_ ( .A(\RegFile/reg_6 [29] ), .Z(\RegFile/_3687_ ) );
BUF_X1 \RegFile/_8885_ ( .A(\RegFile/reg_5 [29] ), .Z(\RegFile/_3655_ ) );
BUF_X1 \RegFile/_8886_ ( .A(\RegFile/reg_4 [29] ), .Z(\RegFile/_3623_ ) );
BUF_X1 \RegFile/_8887_ ( .A(\RegFile/reg_3 [29] ), .Z(\RegFile/_3591_ ) );
BUF_X1 \RegFile/_8888_ ( .A(\RegFile/reg_2 [29] ), .Z(\RegFile/_3559_ ) );
BUF_X1 \RegFile/_8889_ ( .A(\RegFile/reg_1 [29] ), .Z(\RegFile/_3527_ ) );
BUF_X1 \RegFile/_8890_ ( .A(\RegFile/reg_0 [29] ), .Z(\RegFile/_3303_ ) );
BUF_X1 \RegFile/_8891_ ( .A(\RegFile/_0040_ ), .Z(\RegFile/_0104_ ) );
BUF_X1 \RegFile/_8892_ ( .A(\RegFile/_0669_ ), .Z(\_RegFile_io_rd1 [29] ) );
BUF_X1 \RegFile/_8893_ ( .A(\RegFile/_0043_ ), .Z(\RegFile/_0107_ ) );
BUF_X1 \RegFile/_8894_ ( .A(\RegFile/reg_13 [30] ), .Z(\RegFile/_3433_ ) );
BUF_X1 \RegFile/_8895_ ( .A(\RegFile/reg_12 [30] ), .Z(\RegFile/_3401_ ) );
BUF_X1 \RegFile/_8896_ ( .A(\RegFile/reg_11 [30] ), .Z(\RegFile/_3369_ ) );
BUF_X1 \RegFile/_8897_ ( .A(\RegFile/reg_10 [30] ), .Z(\RegFile/_3337_ ) );
BUF_X1 \RegFile/_8898_ ( .A(\RegFile/reg_9 [30] ), .Z(\RegFile/_3785_ ) );
BUF_X1 \RegFile/_8899_ ( .A(\RegFile/reg_8 [30] ), .Z(\RegFile/_3753_ ) );
BUF_X1 \RegFile/_8900_ ( .A(\RegFile/reg_7 [30] ), .Z(\RegFile/_3721_ ) );
BUF_X1 \RegFile/_8901_ ( .A(\RegFile/reg_6 [30] ), .Z(\RegFile/_3689_ ) );
BUF_X1 \RegFile/_8902_ ( .A(\RegFile/reg_5 [30] ), .Z(\RegFile/_3657_ ) );
BUF_X1 \RegFile/_8903_ ( .A(\RegFile/reg_4 [30] ), .Z(\RegFile/_3625_ ) );
BUF_X1 \RegFile/_8904_ ( .A(\RegFile/reg_3 [30] ), .Z(\RegFile/_3593_ ) );
BUF_X1 \RegFile/_8905_ ( .A(\RegFile/reg_2 [30] ), .Z(\RegFile/_3561_ ) );
BUF_X1 \RegFile/_8906_ ( .A(\RegFile/reg_1 [30] ), .Z(\RegFile/_3529_ ) );
BUF_X1 \RegFile/_8907_ ( .A(\RegFile/reg_0 [30] ), .Z(\RegFile/_3305_ ) );
BUF_X1 \RegFile/_8908_ ( .A(\RegFile/_0042_ ), .Z(\RegFile/_0106_ ) );
BUF_X1 \RegFile/_8909_ ( .A(\RegFile/_0671_ ), .Z(\_RegFile_io_rd1 [30] ) );
BUF_X1 \RegFile/_8910_ ( .A(\RegFile/_0045_ ), .Z(\RegFile/_0109_ ) );
BUF_X1 \RegFile/_8911_ ( .A(\RegFile/reg_13 [31] ), .Z(\RegFile/_3434_ ) );
BUF_X1 \RegFile/_8912_ ( .A(\RegFile/reg_12 [31] ), .Z(\RegFile/_3402_ ) );
BUF_X1 \RegFile/_8913_ ( .A(\RegFile/reg_11 [31] ), .Z(\RegFile/_3370_ ) );
BUF_X1 \RegFile/_8914_ ( .A(\RegFile/reg_10 [31] ), .Z(\RegFile/_3338_ ) );
BUF_X1 \RegFile/_8915_ ( .A(\RegFile/reg_9 [31] ), .Z(\RegFile/_3786_ ) );
BUF_X1 \RegFile/_8916_ ( .A(\RegFile/reg_8 [31] ), .Z(\RegFile/_3754_ ) );
BUF_X1 \RegFile/_8917_ ( .A(\RegFile/reg_7 [31] ), .Z(\RegFile/_3722_ ) );
BUF_X1 \RegFile/_8918_ ( .A(\RegFile/reg_6 [31] ), .Z(\RegFile/_3690_ ) );
BUF_X1 \RegFile/_8919_ ( .A(\RegFile/reg_5 [31] ), .Z(\RegFile/_3658_ ) );
BUF_X1 \RegFile/_8920_ ( .A(\RegFile/reg_4 [31] ), .Z(\RegFile/_3626_ ) );
BUF_X1 \RegFile/_8921_ ( .A(\RegFile/reg_3 [31] ), .Z(\RegFile/_3594_ ) );
BUF_X1 \RegFile/_8922_ ( .A(\RegFile/reg_2 [31] ), .Z(\RegFile/_3562_ ) );
BUF_X1 \RegFile/_8923_ ( .A(\RegFile/reg_1 [31] ), .Z(\RegFile/_3530_ ) );
BUF_X1 \RegFile/_8924_ ( .A(\RegFile/reg_0 [31] ), .Z(\RegFile/_3306_ ) );
BUF_X1 \RegFile/_8925_ ( .A(\RegFile/_0044_ ), .Z(\RegFile/_0108_ ) );
BUF_X1 \RegFile/_8926_ ( .A(\RegFile/_0672_ ), .Z(\_RegFile_io_rd1 [31] ) );
BUF_X1 \RegFile/_8927_ ( .A(\_IDU_io_RegFileAccess_ra2 [1] ), .Z(\RegFile/_0645_ ) );
BUF_X1 \RegFile/_8928_ ( .A(\_IDU_io_RegFileAccess_ra2 [0] ), .Z(\RegFile/_0644_ ) );
BUF_X1 \RegFile/_8929_ ( .A(\_IDU_io_RegFileAccess_ra2 [2] ), .Z(\RegFile/_0646_ ) );
BUF_X1 \RegFile/_8930_ ( .A(\_IDU_io_RegFileAccess_ra2 [3] ), .Z(\RegFile/_0647_ ) );
BUF_X1 \RegFile/_8931_ ( .A(\RegFile/_0680_ ), .Z(\_RegFile_io_rd2 [0] ) );
BUF_X1 \RegFile/_8932_ ( .A(\RegFile/_0691_ ), .Z(\_RegFile_io_rd2 [1] ) );
BUF_X1 \RegFile/_8933_ ( .A(\RegFile/_0702_ ), .Z(\_RegFile_io_rd2 [2] ) );
BUF_X1 \RegFile/_8934_ ( .A(\RegFile/_0705_ ), .Z(\_RegFile_io_rd2 [3] ) );
BUF_X1 \RegFile/_8935_ ( .A(\RegFile/_0706_ ), .Z(\_RegFile_io_rd2 [4] ) );
BUF_X1 \RegFile/_8936_ ( .A(\RegFile/_0707_ ), .Z(\_RegFile_io_rd2 [5] ) );
BUF_X1 \RegFile/_8937_ ( .A(\RegFile/_0708_ ), .Z(\_RegFile_io_rd2 [6] ) );
BUF_X1 \RegFile/_8938_ ( .A(\RegFile/_0709_ ), .Z(\_RegFile_io_rd2 [7] ) );
BUF_X1 \RegFile/_8939_ ( .A(\RegFile/_0710_ ), .Z(\_RegFile_io_rd2 [8] ) );
BUF_X1 \RegFile/_8940_ ( .A(\RegFile/_0711_ ), .Z(\_RegFile_io_rd2 [9] ) );
BUF_X1 \RegFile/_8941_ ( .A(\RegFile/_0681_ ), .Z(\_RegFile_io_rd2 [10] ) );
BUF_X1 \RegFile/_8942_ ( .A(\RegFile/_0682_ ), .Z(\_RegFile_io_rd2 [11] ) );
BUF_X1 \RegFile/_8943_ ( .A(\RegFile/_0683_ ), .Z(\_RegFile_io_rd2 [12] ) );
BUF_X1 \RegFile/_8944_ ( .A(\RegFile/_0684_ ), .Z(\_RegFile_io_rd2 [13] ) );
BUF_X1 \RegFile/_8945_ ( .A(\RegFile/_0685_ ), .Z(\_RegFile_io_rd2 [14] ) );
BUF_X1 \RegFile/_8946_ ( .A(\RegFile/_0686_ ), .Z(\_RegFile_io_rd2 [15] ) );
BUF_X1 \RegFile/_8947_ ( .A(\RegFile/_0687_ ), .Z(\_RegFile_io_rd2 [16] ) );
BUF_X1 \RegFile/_8948_ ( .A(\RegFile/_0688_ ), .Z(\_RegFile_io_rd2 [17] ) );
BUF_X1 \RegFile/_8949_ ( .A(\RegFile/_0689_ ), .Z(\_RegFile_io_rd2 [18] ) );
BUF_X1 \RegFile/_8950_ ( .A(\RegFile/_0690_ ), .Z(\_RegFile_io_rd2 [19] ) );
BUF_X1 \RegFile/_8951_ ( .A(\RegFile/_0692_ ), .Z(\_RegFile_io_rd2 [20] ) );
BUF_X1 \RegFile/_8952_ ( .A(\RegFile/_0693_ ), .Z(\_RegFile_io_rd2 [21] ) );
BUF_X1 \RegFile/_8953_ ( .A(\RegFile/_0694_ ), .Z(\_RegFile_io_rd2 [22] ) );
BUF_X1 \RegFile/_8954_ ( .A(\RegFile/_0695_ ), .Z(\_RegFile_io_rd2 [23] ) );
BUF_X1 \RegFile/_8955_ ( .A(\RegFile/_0696_ ), .Z(\_RegFile_io_rd2 [24] ) );
BUF_X1 \RegFile/_8956_ ( .A(\RegFile/_0697_ ), .Z(\_RegFile_io_rd2 [25] ) );
BUF_X1 \RegFile/_8957_ ( .A(\RegFile/_0698_ ), .Z(\_RegFile_io_rd2 [26] ) );
BUF_X1 \RegFile/_8958_ ( .A(\RegFile/_0699_ ), .Z(\_RegFile_io_rd2 [27] ) );
BUF_X1 \RegFile/_8959_ ( .A(\RegFile/_0700_ ), .Z(\_RegFile_io_rd2 [28] ) );
BUF_X1 \RegFile/_8960_ ( .A(\RegFile/_0701_ ), .Z(\_RegFile_io_rd2 [29] ) );
BUF_X1 \RegFile/_8961_ ( .A(\RegFile/_0703_ ), .Z(\_RegFile_io_rd2 [30] ) );
BUF_X1 \RegFile/_8962_ ( .A(\RegFile/_0704_ ), .Z(\_RegFile_io_rd2 [31] ) );
BUF_X1 \RegFile/_8963_ ( .A(\RegFile/reg_14 [0] ), .Z(\RegFile/_3442_ ) );
BUF_X1 \RegFile/_8964_ ( .A(\RegFile/reg_15 [0] ), .Z(\RegFile/_3474_ ) );
BUF_X1 \RegFile/_8965_ ( .A(_WBU_io_RegFileAccess_we ), .Z(\RegFile/_0748_ ) );
BUF_X1 \RegFile/_8966_ ( .A(\_WBU_io_RegFileAccess_wd [0] ), .Z(\RegFile/_0716_ ) );
BUF_X1 \RegFile/_8967_ ( .A(\RegFile/reg_14 [1] ), .Z(\RegFile/_3453_ ) );
BUF_X1 \RegFile/_8968_ ( .A(\RegFile/reg_15 [1] ), .Z(\RegFile/_3485_ ) );
BUF_X1 \RegFile/_8969_ ( .A(\_WBU_io_RegFileAccess_wd [1] ), .Z(\RegFile/_0727_ ) );
BUF_X1 \RegFile/_8970_ ( .A(\RegFile/reg_14 [2] ), .Z(\RegFile/_3464_ ) );
BUF_X1 \RegFile/_8971_ ( .A(\RegFile/reg_15 [2] ), .Z(\RegFile/_3496_ ) );
BUF_X1 \RegFile/_8972_ ( .A(\_WBU_io_RegFileAccess_wd [2] ), .Z(\RegFile/_0738_ ) );
BUF_X1 \RegFile/_8973_ ( .A(\RegFile/reg_14 [3] ), .Z(\RegFile/_3467_ ) );
BUF_X1 \RegFile/_8974_ ( .A(\RegFile/reg_15 [3] ), .Z(\RegFile/_3499_ ) );
BUF_X1 \RegFile/_8975_ ( .A(\_WBU_io_RegFileAccess_wd [3] ), .Z(\RegFile/_0741_ ) );
BUF_X1 \RegFile/_8976_ ( .A(\RegFile/reg_14 [4] ), .Z(\RegFile/_3468_ ) );
BUF_X1 \RegFile/_8977_ ( .A(\RegFile/reg_15 [4] ), .Z(\RegFile/_3500_ ) );
BUF_X1 \RegFile/_8978_ ( .A(\_WBU_io_RegFileAccess_wd [4] ), .Z(\RegFile/_0742_ ) );
BUF_X1 \RegFile/_8979_ ( .A(\RegFile/reg_14 [5] ), .Z(\RegFile/_3469_ ) );
BUF_X1 \RegFile/_8980_ ( .A(\RegFile/reg_15 [5] ), .Z(\RegFile/_3501_ ) );
BUF_X1 \RegFile/_8981_ ( .A(\_WBU_io_RegFileAccess_wd [5] ), .Z(\RegFile/_0743_ ) );
BUF_X1 \RegFile/_8982_ ( .A(\RegFile/reg_14 [6] ), .Z(\RegFile/_3470_ ) );
BUF_X1 \RegFile/_8983_ ( .A(\RegFile/reg_15 [6] ), .Z(\RegFile/_3502_ ) );
BUF_X1 \RegFile/_8984_ ( .A(\_WBU_io_RegFileAccess_wd [6] ), .Z(\RegFile/_0744_ ) );
BUF_X1 \RegFile/_8985_ ( .A(\RegFile/reg_14 [7] ), .Z(\RegFile/_3471_ ) );
BUF_X1 \RegFile/_8986_ ( .A(\RegFile/reg_15 [7] ), .Z(\RegFile/_3503_ ) );
BUF_X1 \RegFile/_8987_ ( .A(\_WBU_io_RegFileAccess_wd [7] ), .Z(\RegFile/_0745_ ) );
BUF_X1 \RegFile/_8988_ ( .A(\RegFile/reg_14 [8] ), .Z(\RegFile/_3472_ ) );
BUF_X1 \RegFile/_8989_ ( .A(\RegFile/reg_15 [8] ), .Z(\RegFile/_3504_ ) );
BUF_X1 \RegFile/_8990_ ( .A(\_WBU_io_RegFileAccess_wd [8] ), .Z(\RegFile/_0746_ ) );
BUF_X1 \RegFile/_8991_ ( .A(\RegFile/reg_14 [9] ), .Z(\RegFile/_3473_ ) );
BUF_X1 \RegFile/_8992_ ( .A(\RegFile/reg_15 [9] ), .Z(\RegFile/_3505_ ) );
BUF_X1 \RegFile/_8993_ ( .A(\_WBU_io_RegFileAccess_wd [9] ), .Z(\RegFile/_0747_ ) );
BUF_X1 \RegFile/_8994_ ( .A(\RegFile/reg_14 [10] ), .Z(\RegFile/_3443_ ) );
BUF_X1 \RegFile/_8995_ ( .A(\RegFile/reg_15 [10] ), .Z(\RegFile/_3475_ ) );
BUF_X1 \RegFile/_8996_ ( .A(\_WBU_io_RegFileAccess_wd [10] ), .Z(\RegFile/_0717_ ) );
BUF_X1 \RegFile/_8997_ ( .A(\RegFile/reg_14 [11] ), .Z(\RegFile/_3444_ ) );
BUF_X1 \RegFile/_8998_ ( .A(\RegFile/reg_15 [11] ), .Z(\RegFile/_3476_ ) );
BUF_X1 \RegFile/_8999_ ( .A(\_WBU_io_RegFileAccess_wd [11] ), .Z(\RegFile/_0718_ ) );
BUF_X1 \RegFile/_9000_ ( .A(\RegFile/reg_14 [12] ), .Z(\RegFile/_3445_ ) );
BUF_X1 \RegFile/_9001_ ( .A(\RegFile/reg_15 [12] ), .Z(\RegFile/_3477_ ) );
BUF_X1 \RegFile/_9002_ ( .A(\_WBU_io_RegFileAccess_wd [12] ), .Z(\RegFile/_0719_ ) );
BUF_X1 \RegFile/_9003_ ( .A(\RegFile/reg_14 [13] ), .Z(\RegFile/_3446_ ) );
BUF_X1 \RegFile/_9004_ ( .A(\RegFile/reg_15 [13] ), .Z(\RegFile/_3478_ ) );
BUF_X1 \RegFile/_9005_ ( .A(\_WBU_io_RegFileAccess_wd [13] ), .Z(\RegFile/_0720_ ) );
BUF_X1 \RegFile/_9006_ ( .A(\RegFile/reg_14 [14] ), .Z(\RegFile/_3447_ ) );
BUF_X1 \RegFile/_9007_ ( .A(\RegFile/reg_15 [14] ), .Z(\RegFile/_3479_ ) );
BUF_X1 \RegFile/_9008_ ( .A(\_WBU_io_RegFileAccess_wd [14] ), .Z(\RegFile/_0721_ ) );
BUF_X1 \RegFile/_9009_ ( .A(\RegFile/reg_14 [15] ), .Z(\RegFile/_3448_ ) );
BUF_X1 \RegFile/_9010_ ( .A(\RegFile/reg_15 [15] ), .Z(\RegFile/_3480_ ) );
BUF_X1 \RegFile/_9011_ ( .A(\_WBU_io_RegFileAccess_wd [15] ), .Z(\RegFile/_0722_ ) );
BUF_X1 \RegFile/_9012_ ( .A(\RegFile/reg_14 [16] ), .Z(\RegFile/_3449_ ) );
BUF_X1 \RegFile/_9013_ ( .A(\RegFile/reg_15 [16] ), .Z(\RegFile/_3481_ ) );
BUF_X1 \RegFile/_9014_ ( .A(\_WBU_io_RegFileAccess_wd [16] ), .Z(\RegFile/_0723_ ) );
BUF_X1 \RegFile/_9015_ ( .A(\RegFile/reg_14 [17] ), .Z(\RegFile/_3450_ ) );
BUF_X1 \RegFile/_9016_ ( .A(\RegFile/reg_15 [17] ), .Z(\RegFile/_3482_ ) );
BUF_X1 \RegFile/_9017_ ( .A(\_WBU_io_RegFileAccess_wd [17] ), .Z(\RegFile/_0724_ ) );
BUF_X1 \RegFile/_9018_ ( .A(\RegFile/reg_14 [18] ), .Z(\RegFile/_3451_ ) );
BUF_X1 \RegFile/_9019_ ( .A(\RegFile/reg_15 [18] ), .Z(\RegFile/_3483_ ) );
BUF_X1 \RegFile/_9020_ ( .A(\_WBU_io_RegFileAccess_wd [18] ), .Z(\RegFile/_0725_ ) );
BUF_X1 \RegFile/_9021_ ( .A(\RegFile/reg_14 [19] ), .Z(\RegFile/_3452_ ) );
BUF_X1 \RegFile/_9022_ ( .A(\RegFile/reg_15 [19] ), .Z(\RegFile/_3484_ ) );
BUF_X1 \RegFile/_9023_ ( .A(\_WBU_io_RegFileAccess_wd [19] ), .Z(\RegFile/_0726_ ) );
BUF_X1 \RegFile/_9024_ ( .A(\RegFile/reg_14 [20] ), .Z(\RegFile/_3454_ ) );
BUF_X1 \RegFile/_9025_ ( .A(\RegFile/reg_15 [20] ), .Z(\RegFile/_3486_ ) );
BUF_X1 \RegFile/_9026_ ( .A(\_WBU_io_RegFileAccess_wd [20] ), .Z(\RegFile/_0728_ ) );
BUF_X1 \RegFile/_9027_ ( .A(\RegFile/reg_14 [21] ), .Z(\RegFile/_3455_ ) );
BUF_X1 \RegFile/_9028_ ( .A(\RegFile/reg_15 [21] ), .Z(\RegFile/_3487_ ) );
BUF_X1 \RegFile/_9029_ ( .A(\_WBU_io_RegFileAccess_wd [21] ), .Z(\RegFile/_0729_ ) );
BUF_X1 \RegFile/_9030_ ( .A(\RegFile/reg_14 [22] ), .Z(\RegFile/_3456_ ) );
BUF_X1 \RegFile/_9031_ ( .A(\RegFile/reg_15 [22] ), .Z(\RegFile/_3488_ ) );
BUF_X1 \RegFile/_9032_ ( .A(\_WBU_io_RegFileAccess_wd [22] ), .Z(\RegFile/_0730_ ) );
BUF_X1 \RegFile/_9033_ ( .A(\RegFile/reg_14 [23] ), .Z(\RegFile/_3457_ ) );
BUF_X1 \RegFile/_9034_ ( .A(\RegFile/reg_15 [23] ), .Z(\RegFile/_3489_ ) );
BUF_X1 \RegFile/_9035_ ( .A(\_WBU_io_RegFileAccess_wd [23] ), .Z(\RegFile/_0731_ ) );
BUF_X1 \RegFile/_9036_ ( .A(\RegFile/reg_14 [24] ), .Z(\RegFile/_3458_ ) );
BUF_X1 \RegFile/_9037_ ( .A(\RegFile/reg_15 [24] ), .Z(\RegFile/_3490_ ) );
BUF_X1 \RegFile/_9038_ ( .A(\_WBU_io_RegFileAccess_wd [24] ), .Z(\RegFile/_0732_ ) );
BUF_X1 \RegFile/_9039_ ( .A(\RegFile/reg_14 [25] ), .Z(\RegFile/_3459_ ) );
BUF_X1 \RegFile/_9040_ ( .A(\RegFile/reg_15 [25] ), .Z(\RegFile/_3491_ ) );
BUF_X1 \RegFile/_9041_ ( .A(\_WBU_io_RegFileAccess_wd [25] ), .Z(\RegFile/_0733_ ) );
BUF_X1 \RegFile/_9042_ ( .A(\RegFile/reg_14 [26] ), .Z(\RegFile/_3460_ ) );
BUF_X1 \RegFile/_9043_ ( .A(\RegFile/reg_15 [26] ), .Z(\RegFile/_3492_ ) );
BUF_X1 \RegFile/_9044_ ( .A(\_WBU_io_RegFileAccess_wd [26] ), .Z(\RegFile/_0734_ ) );
BUF_X1 \RegFile/_9045_ ( .A(\RegFile/reg_14 [27] ), .Z(\RegFile/_3461_ ) );
BUF_X1 \RegFile/_9046_ ( .A(\RegFile/reg_15 [27] ), .Z(\RegFile/_3493_ ) );
BUF_X1 \RegFile/_9047_ ( .A(\_WBU_io_RegFileAccess_wd [27] ), .Z(\RegFile/_0735_ ) );
BUF_X1 \RegFile/_9048_ ( .A(\RegFile/reg_14 [28] ), .Z(\RegFile/_3462_ ) );
BUF_X1 \RegFile/_9049_ ( .A(\RegFile/reg_15 [28] ), .Z(\RegFile/_3494_ ) );
BUF_X1 \RegFile/_9050_ ( .A(\_WBU_io_RegFileAccess_wd [28] ), .Z(\RegFile/_0736_ ) );
BUF_X1 \RegFile/_9051_ ( .A(\RegFile/reg_14 [29] ), .Z(\RegFile/_3463_ ) );
BUF_X1 \RegFile/_9052_ ( .A(\RegFile/reg_15 [29] ), .Z(\RegFile/_3495_ ) );
BUF_X1 \RegFile/_9053_ ( .A(\_WBU_io_RegFileAccess_wd [29] ), .Z(\RegFile/_0737_ ) );
BUF_X1 \RegFile/_9054_ ( .A(\RegFile/reg_14 [30] ), .Z(\RegFile/_3465_ ) );
BUF_X1 \RegFile/_9055_ ( .A(\RegFile/reg_15 [30] ), .Z(\RegFile/_3497_ ) );
BUF_X1 \RegFile/_9056_ ( .A(\_WBU_io_RegFileAccess_wd [30] ), .Z(\RegFile/_0739_ ) );
BUF_X1 \RegFile/_9057_ ( .A(\RegFile/reg_14 [31] ), .Z(\RegFile/_3466_ ) );
BUF_X1 \RegFile/_9058_ ( .A(\RegFile/reg_15 [31] ), .Z(\RegFile/_3498_ ) );
BUF_X1 \RegFile/_9059_ ( .A(\_WBU_io_RegFileAccess_wd [31] ), .Z(\RegFile/_0740_ ) );
BUF_X1 \RegFile/_9060_ ( .A(\RegFile/_0608_ ), .Z(\RegFile/_4722_ ) );
BUF_X1 \RegFile/_9061_ ( .A(\RegFile/_0609_ ), .Z(\RegFile/_4723_ ) );
BUF_X1 \RegFile/_9062_ ( .A(\RegFile/_0610_ ), .Z(\RegFile/_4724_ ) );
BUF_X1 \RegFile/_9063_ ( .A(\RegFile/_0611_ ), .Z(\RegFile/_4725_ ) );
BUF_X1 \RegFile/_9064_ ( .A(\RegFile/_0612_ ), .Z(\RegFile/_4726_ ) );
BUF_X1 \RegFile/_9065_ ( .A(\RegFile/_0613_ ), .Z(\RegFile/_4727_ ) );
BUF_X1 \RegFile/_9066_ ( .A(\RegFile/_0614_ ), .Z(\RegFile/_4728_ ) );
BUF_X1 \RegFile/_9067_ ( .A(\RegFile/_0615_ ), .Z(\RegFile/_4729_ ) );
BUF_X1 \RegFile/_9068_ ( .A(\RegFile/_0616_ ), .Z(\RegFile/_4730_ ) );
BUF_X1 \RegFile/_9069_ ( .A(\RegFile/_0617_ ), .Z(\RegFile/_4731_ ) );
BUF_X1 \RegFile/_9070_ ( .A(\RegFile/_0618_ ), .Z(\RegFile/_4732_ ) );
BUF_X1 \RegFile/_9071_ ( .A(\RegFile/_0619_ ), .Z(\RegFile/_4733_ ) );
BUF_X1 \RegFile/_9072_ ( .A(\RegFile/_0620_ ), .Z(\RegFile/_4734_ ) );
BUF_X1 \RegFile/_9073_ ( .A(\RegFile/_0621_ ), .Z(\RegFile/_4735_ ) );
BUF_X1 \RegFile/_9074_ ( .A(\RegFile/_0622_ ), .Z(\RegFile/_4736_ ) );
BUF_X1 \RegFile/_9075_ ( .A(\RegFile/_0623_ ), .Z(\RegFile/_4737_ ) );
BUF_X1 \RegFile/_9076_ ( .A(\RegFile/_0624_ ), .Z(\RegFile/_4738_ ) );
BUF_X1 \RegFile/_9077_ ( .A(\RegFile/_0625_ ), .Z(\RegFile/_4739_ ) );
BUF_X1 \RegFile/_9078_ ( .A(\RegFile/_0626_ ), .Z(\RegFile/_4740_ ) );
BUF_X1 \RegFile/_9079_ ( .A(\RegFile/_0627_ ), .Z(\RegFile/_4741_ ) );
BUF_X1 \RegFile/_9080_ ( .A(\RegFile/_0628_ ), .Z(\RegFile/_4742_ ) );
BUF_X1 \RegFile/_9081_ ( .A(\RegFile/_0629_ ), .Z(\RegFile/_4743_ ) );
BUF_X1 \RegFile/_9082_ ( .A(\RegFile/_0630_ ), .Z(\RegFile/_4744_ ) );
BUF_X1 \RegFile/_9083_ ( .A(\RegFile/_0631_ ), .Z(\RegFile/_4745_ ) );
BUF_X1 \RegFile/_9084_ ( .A(\RegFile/_0632_ ), .Z(\RegFile/_4746_ ) );
BUF_X1 \RegFile/_9085_ ( .A(\RegFile/_0633_ ), .Z(\RegFile/_4747_ ) );
BUF_X1 \RegFile/_9086_ ( .A(\RegFile/_0634_ ), .Z(\RegFile/_4748_ ) );
BUF_X1 \RegFile/_9087_ ( .A(\RegFile/_0635_ ), .Z(\RegFile/_4749_ ) );
BUF_X1 \RegFile/_9088_ ( .A(\RegFile/_0636_ ), .Z(\RegFile/_4750_ ) );
BUF_X1 \RegFile/_9089_ ( .A(\RegFile/_0637_ ), .Z(\RegFile/_4751_ ) );
BUF_X1 \RegFile/_9090_ ( .A(\RegFile/_0638_ ), .Z(\RegFile/_4752_ ) );
BUF_X1 \RegFile/_9091_ ( .A(\RegFile/_0639_ ), .Z(\RegFile/_4753_ ) );
BUF_X1 \RegFile/_9092_ ( .A(\RegFile/_0128_ ), .Z(\RegFile/_4242_ ) );
BUF_X1 \RegFile/_9093_ ( .A(\RegFile/_0129_ ), .Z(\RegFile/_4243_ ) );
BUF_X1 \RegFile/_9094_ ( .A(\RegFile/_0130_ ), .Z(\RegFile/_4244_ ) );
BUF_X1 \RegFile/_9095_ ( .A(\RegFile/_0131_ ), .Z(\RegFile/_4245_ ) );
BUF_X1 \RegFile/_9096_ ( .A(\RegFile/_0132_ ), .Z(\RegFile/_4246_ ) );
BUF_X1 \RegFile/_9097_ ( .A(\RegFile/_0133_ ), .Z(\RegFile/_4247_ ) );
BUF_X1 \RegFile/_9098_ ( .A(\RegFile/_0134_ ), .Z(\RegFile/_4248_ ) );
BUF_X1 \RegFile/_9099_ ( .A(\RegFile/_0135_ ), .Z(\RegFile/_4249_ ) );
BUF_X1 \RegFile/_9100_ ( .A(\RegFile/_0136_ ), .Z(\RegFile/_4250_ ) );
BUF_X1 \RegFile/_9101_ ( .A(\RegFile/_0137_ ), .Z(\RegFile/_4251_ ) );
BUF_X1 \RegFile/_9102_ ( .A(\RegFile/_0138_ ), .Z(\RegFile/_4252_ ) );
BUF_X1 \RegFile/_9103_ ( .A(\RegFile/_0139_ ), .Z(\RegFile/_4253_ ) );
BUF_X1 \RegFile/_9104_ ( .A(\RegFile/_0140_ ), .Z(\RegFile/_4254_ ) );
BUF_X1 \RegFile/_9105_ ( .A(\RegFile/_0141_ ), .Z(\RegFile/_4255_ ) );
BUF_X1 \RegFile/_9106_ ( .A(\RegFile/_0142_ ), .Z(\RegFile/_4256_ ) );
BUF_X1 \RegFile/_9107_ ( .A(\RegFile/_0143_ ), .Z(\RegFile/_4257_ ) );
BUF_X1 \RegFile/_9108_ ( .A(\RegFile/_0144_ ), .Z(\RegFile/_4258_ ) );
BUF_X1 \RegFile/_9109_ ( .A(\RegFile/_0145_ ), .Z(\RegFile/_4259_ ) );
BUF_X1 \RegFile/_9110_ ( .A(\RegFile/_0146_ ), .Z(\RegFile/_4260_ ) );
BUF_X1 \RegFile/_9111_ ( .A(\RegFile/_0147_ ), .Z(\RegFile/_4261_ ) );
BUF_X1 \RegFile/_9112_ ( .A(\RegFile/_0148_ ), .Z(\RegFile/_4262_ ) );
BUF_X1 \RegFile/_9113_ ( .A(\RegFile/_0149_ ), .Z(\RegFile/_4263_ ) );
BUF_X1 \RegFile/_9114_ ( .A(\RegFile/_0150_ ), .Z(\RegFile/_4264_ ) );
BUF_X1 \RegFile/_9115_ ( .A(\RegFile/_0151_ ), .Z(\RegFile/_4265_ ) );
BUF_X1 \RegFile/_9116_ ( .A(\RegFile/_0152_ ), .Z(\RegFile/_4266_ ) );
BUF_X1 \RegFile/_9117_ ( .A(\RegFile/_0153_ ), .Z(\RegFile/_4267_ ) );
BUF_X1 \RegFile/_9118_ ( .A(\RegFile/_0154_ ), .Z(\RegFile/_4268_ ) );
BUF_X1 \RegFile/_9119_ ( .A(\RegFile/_0155_ ), .Z(\RegFile/_4269_ ) );
BUF_X1 \RegFile/_9120_ ( .A(\RegFile/_0156_ ), .Z(\RegFile/_4270_ ) );
BUF_X1 \RegFile/_9121_ ( .A(\RegFile/_0157_ ), .Z(\RegFile/_4271_ ) );
BUF_X1 \RegFile/_9122_ ( .A(\RegFile/_0158_ ), .Z(\RegFile/_4272_ ) );
BUF_X1 \RegFile/_9123_ ( .A(\RegFile/_0159_ ), .Z(\RegFile/_4273_ ) );
BUF_X1 \RegFile/_9124_ ( .A(\RegFile/_0160_ ), .Z(\RegFile/_4274_ ) );
BUF_X1 \RegFile/_9125_ ( .A(\RegFile/_0161_ ), .Z(\RegFile/_4275_ ) );
BUF_X1 \RegFile/_9126_ ( .A(\RegFile/_0162_ ), .Z(\RegFile/_4276_ ) );
BUF_X1 \RegFile/_9127_ ( .A(\RegFile/_0163_ ), .Z(\RegFile/_4277_ ) );
BUF_X1 \RegFile/_9128_ ( .A(\RegFile/_0164_ ), .Z(\RegFile/_4278_ ) );
BUF_X1 \RegFile/_9129_ ( .A(\RegFile/_0165_ ), .Z(\RegFile/_4279_ ) );
BUF_X1 \RegFile/_9130_ ( .A(\RegFile/_0166_ ), .Z(\RegFile/_4280_ ) );
BUF_X1 \RegFile/_9131_ ( .A(\RegFile/_0167_ ), .Z(\RegFile/_4281_ ) );
BUF_X1 \RegFile/_9132_ ( .A(\RegFile/_0168_ ), .Z(\RegFile/_4282_ ) );
BUF_X1 \RegFile/_9133_ ( .A(\RegFile/_0169_ ), .Z(\RegFile/_4283_ ) );
BUF_X1 \RegFile/_9134_ ( .A(\RegFile/_0170_ ), .Z(\RegFile/_4284_ ) );
BUF_X1 \RegFile/_9135_ ( .A(\RegFile/_0171_ ), .Z(\RegFile/_4285_ ) );
BUF_X1 \RegFile/_9136_ ( .A(\RegFile/_0172_ ), .Z(\RegFile/_4286_ ) );
BUF_X1 \RegFile/_9137_ ( .A(\RegFile/_0173_ ), .Z(\RegFile/_4287_ ) );
BUF_X1 \RegFile/_9138_ ( .A(\RegFile/_0174_ ), .Z(\RegFile/_4288_ ) );
BUF_X1 \RegFile/_9139_ ( .A(\RegFile/_0175_ ), .Z(\RegFile/_4289_ ) );
BUF_X1 \RegFile/_9140_ ( .A(\RegFile/_0176_ ), .Z(\RegFile/_4290_ ) );
BUF_X1 \RegFile/_9141_ ( .A(\RegFile/_0177_ ), .Z(\RegFile/_4291_ ) );
BUF_X1 \RegFile/_9142_ ( .A(\RegFile/_0178_ ), .Z(\RegFile/_4292_ ) );
BUF_X1 \RegFile/_9143_ ( .A(\RegFile/_0179_ ), .Z(\RegFile/_4293_ ) );
BUF_X1 \RegFile/_9144_ ( .A(\RegFile/_0180_ ), .Z(\RegFile/_4294_ ) );
BUF_X1 \RegFile/_9145_ ( .A(\RegFile/_0181_ ), .Z(\RegFile/_4295_ ) );
BUF_X1 \RegFile/_9146_ ( .A(\RegFile/_0182_ ), .Z(\RegFile/_4296_ ) );
BUF_X1 \RegFile/_9147_ ( .A(\RegFile/_0183_ ), .Z(\RegFile/_4297_ ) );
BUF_X1 \RegFile/_9148_ ( .A(\RegFile/_0184_ ), .Z(\RegFile/_4298_ ) );
BUF_X1 \RegFile/_9149_ ( .A(\RegFile/_0185_ ), .Z(\RegFile/_4299_ ) );
BUF_X1 \RegFile/_9150_ ( .A(\RegFile/_0186_ ), .Z(\RegFile/_4300_ ) );
BUF_X1 \RegFile/_9151_ ( .A(\RegFile/_0187_ ), .Z(\RegFile/_4301_ ) );
BUF_X1 \RegFile/_9152_ ( .A(\RegFile/_0188_ ), .Z(\RegFile/_4302_ ) );
BUF_X1 \RegFile/_9153_ ( .A(\RegFile/_0189_ ), .Z(\RegFile/_4303_ ) );
BUF_X1 \RegFile/_9154_ ( .A(\RegFile/_0190_ ), .Z(\RegFile/_4304_ ) );
BUF_X1 \RegFile/_9155_ ( .A(\RegFile/_0191_ ), .Z(\RegFile/_4305_ ) );
BUF_X1 \RegFile/_9156_ ( .A(\RegFile/_0192_ ), .Z(\RegFile/_4306_ ) );
BUF_X1 \RegFile/_9157_ ( .A(\RegFile/_0193_ ), .Z(\RegFile/_4307_ ) );
BUF_X1 \RegFile/_9158_ ( .A(\RegFile/_0194_ ), .Z(\RegFile/_4308_ ) );
BUF_X1 \RegFile/_9159_ ( .A(\RegFile/_0195_ ), .Z(\RegFile/_4309_ ) );
BUF_X1 \RegFile/_9160_ ( .A(\RegFile/_0196_ ), .Z(\RegFile/_4310_ ) );
BUF_X1 \RegFile/_9161_ ( .A(\RegFile/_0197_ ), .Z(\RegFile/_4311_ ) );
BUF_X1 \RegFile/_9162_ ( .A(\RegFile/_0198_ ), .Z(\RegFile/_4312_ ) );
BUF_X1 \RegFile/_9163_ ( .A(\RegFile/_0199_ ), .Z(\RegFile/_4313_ ) );
BUF_X1 \RegFile/_9164_ ( .A(\RegFile/_0200_ ), .Z(\RegFile/_4314_ ) );
BUF_X1 \RegFile/_9165_ ( .A(\RegFile/_0201_ ), .Z(\RegFile/_4315_ ) );
BUF_X1 \RegFile/_9166_ ( .A(\RegFile/_0202_ ), .Z(\RegFile/_4316_ ) );
BUF_X1 \RegFile/_9167_ ( .A(\RegFile/_0203_ ), .Z(\RegFile/_4317_ ) );
BUF_X1 \RegFile/_9168_ ( .A(\RegFile/_0204_ ), .Z(\RegFile/_4318_ ) );
BUF_X1 \RegFile/_9169_ ( .A(\RegFile/_0205_ ), .Z(\RegFile/_4319_ ) );
BUF_X1 \RegFile/_9170_ ( .A(\RegFile/_0206_ ), .Z(\RegFile/_4320_ ) );
BUF_X1 \RegFile/_9171_ ( .A(\RegFile/_0207_ ), .Z(\RegFile/_4321_ ) );
BUF_X1 \RegFile/_9172_ ( .A(\RegFile/_0208_ ), .Z(\RegFile/_4322_ ) );
BUF_X1 \RegFile/_9173_ ( .A(\RegFile/_0209_ ), .Z(\RegFile/_4323_ ) );
BUF_X1 \RegFile/_9174_ ( .A(\RegFile/_0210_ ), .Z(\RegFile/_4324_ ) );
BUF_X1 \RegFile/_9175_ ( .A(\RegFile/_0211_ ), .Z(\RegFile/_4325_ ) );
BUF_X1 \RegFile/_9176_ ( .A(\RegFile/_0212_ ), .Z(\RegFile/_4326_ ) );
BUF_X1 \RegFile/_9177_ ( .A(\RegFile/_0213_ ), .Z(\RegFile/_4327_ ) );
BUF_X1 \RegFile/_9178_ ( .A(\RegFile/_0214_ ), .Z(\RegFile/_4328_ ) );
BUF_X1 \RegFile/_9179_ ( .A(\RegFile/_0215_ ), .Z(\RegFile/_4329_ ) );
BUF_X1 \RegFile/_9180_ ( .A(\RegFile/_0216_ ), .Z(\RegFile/_4330_ ) );
BUF_X1 \RegFile/_9181_ ( .A(\RegFile/_0217_ ), .Z(\RegFile/_4331_ ) );
BUF_X1 \RegFile/_9182_ ( .A(\RegFile/_0218_ ), .Z(\RegFile/_4332_ ) );
BUF_X1 \RegFile/_9183_ ( .A(\RegFile/_0219_ ), .Z(\RegFile/_4333_ ) );
BUF_X1 \RegFile/_9184_ ( .A(\RegFile/_0220_ ), .Z(\RegFile/_4334_ ) );
BUF_X1 \RegFile/_9185_ ( .A(\RegFile/_0221_ ), .Z(\RegFile/_4335_ ) );
BUF_X1 \RegFile/_9186_ ( .A(\RegFile/_0222_ ), .Z(\RegFile/_4336_ ) );
BUF_X1 \RegFile/_9187_ ( .A(\RegFile/_0223_ ), .Z(\RegFile/_4337_ ) );
BUF_X1 \RegFile/_9188_ ( .A(\RegFile/_0224_ ), .Z(\RegFile/_4338_ ) );
BUF_X1 \RegFile/_9189_ ( .A(\RegFile/_0225_ ), .Z(\RegFile/_4339_ ) );
BUF_X1 \RegFile/_9190_ ( .A(\RegFile/_0226_ ), .Z(\RegFile/_4340_ ) );
BUF_X1 \RegFile/_9191_ ( .A(\RegFile/_0227_ ), .Z(\RegFile/_4341_ ) );
BUF_X1 \RegFile/_9192_ ( .A(\RegFile/_0228_ ), .Z(\RegFile/_4342_ ) );
BUF_X1 \RegFile/_9193_ ( .A(\RegFile/_0229_ ), .Z(\RegFile/_4343_ ) );
BUF_X1 \RegFile/_9194_ ( .A(\RegFile/_0230_ ), .Z(\RegFile/_4344_ ) );
BUF_X1 \RegFile/_9195_ ( .A(\RegFile/_0231_ ), .Z(\RegFile/_4345_ ) );
BUF_X1 \RegFile/_9196_ ( .A(\RegFile/_0232_ ), .Z(\RegFile/_4346_ ) );
BUF_X1 \RegFile/_9197_ ( .A(\RegFile/_0233_ ), .Z(\RegFile/_4347_ ) );
BUF_X1 \RegFile/_9198_ ( .A(\RegFile/_0234_ ), .Z(\RegFile/_4348_ ) );
BUF_X1 \RegFile/_9199_ ( .A(\RegFile/_0235_ ), .Z(\RegFile/_4349_ ) );
BUF_X1 \RegFile/_9200_ ( .A(\RegFile/_0236_ ), .Z(\RegFile/_4350_ ) );
BUF_X1 \RegFile/_9201_ ( .A(\RegFile/_0237_ ), .Z(\RegFile/_4351_ ) );
BUF_X1 \RegFile/_9202_ ( .A(\RegFile/_0238_ ), .Z(\RegFile/_4352_ ) );
BUF_X1 \RegFile/_9203_ ( .A(\RegFile/_0239_ ), .Z(\RegFile/_4353_ ) );
BUF_X1 \RegFile/_9204_ ( .A(\RegFile/_0240_ ), .Z(\RegFile/_4354_ ) );
BUF_X1 \RegFile/_9205_ ( .A(\RegFile/_0241_ ), .Z(\RegFile/_4355_ ) );
BUF_X1 \RegFile/_9206_ ( .A(\RegFile/_0242_ ), .Z(\RegFile/_4356_ ) );
BUF_X1 \RegFile/_9207_ ( .A(\RegFile/_0243_ ), .Z(\RegFile/_4357_ ) );
BUF_X1 \RegFile/_9208_ ( .A(\RegFile/_0244_ ), .Z(\RegFile/_4358_ ) );
BUF_X1 \RegFile/_9209_ ( .A(\RegFile/_0245_ ), .Z(\RegFile/_4359_ ) );
BUF_X1 \RegFile/_9210_ ( .A(\RegFile/_0246_ ), .Z(\RegFile/_4360_ ) );
BUF_X1 \RegFile/_9211_ ( .A(\RegFile/_0247_ ), .Z(\RegFile/_4361_ ) );
BUF_X1 \RegFile/_9212_ ( .A(\RegFile/_0248_ ), .Z(\RegFile/_4362_ ) );
BUF_X1 \RegFile/_9213_ ( .A(\RegFile/_0249_ ), .Z(\RegFile/_4363_ ) );
BUF_X1 \RegFile/_9214_ ( .A(\RegFile/_0250_ ), .Z(\RegFile/_4364_ ) );
BUF_X1 \RegFile/_9215_ ( .A(\RegFile/_0251_ ), .Z(\RegFile/_4365_ ) );
BUF_X1 \RegFile/_9216_ ( .A(\RegFile/_0252_ ), .Z(\RegFile/_4366_ ) );
BUF_X1 \RegFile/_9217_ ( .A(\RegFile/_0253_ ), .Z(\RegFile/_4367_ ) );
BUF_X1 \RegFile/_9218_ ( .A(\RegFile/_0254_ ), .Z(\RegFile/_4368_ ) );
BUF_X1 \RegFile/_9219_ ( .A(\RegFile/_0255_ ), .Z(\RegFile/_4369_ ) );
BUF_X1 \RegFile/_9220_ ( .A(\RegFile/_0256_ ), .Z(\RegFile/_4370_ ) );
BUF_X1 \RegFile/_9221_ ( .A(\RegFile/_0257_ ), .Z(\RegFile/_4371_ ) );
BUF_X1 \RegFile/_9222_ ( .A(\RegFile/_0258_ ), .Z(\RegFile/_4372_ ) );
BUF_X1 \RegFile/_9223_ ( .A(\RegFile/_0259_ ), .Z(\RegFile/_4373_ ) );
BUF_X1 \RegFile/_9224_ ( .A(\RegFile/_0260_ ), .Z(\RegFile/_4374_ ) );
BUF_X1 \RegFile/_9225_ ( .A(\RegFile/_0261_ ), .Z(\RegFile/_4375_ ) );
BUF_X1 \RegFile/_9226_ ( .A(\RegFile/_0262_ ), .Z(\RegFile/_4376_ ) );
BUF_X1 \RegFile/_9227_ ( .A(\RegFile/_0263_ ), .Z(\RegFile/_4377_ ) );
BUF_X1 \RegFile/_9228_ ( .A(\RegFile/_0264_ ), .Z(\RegFile/_4378_ ) );
BUF_X1 \RegFile/_9229_ ( .A(\RegFile/_0265_ ), .Z(\RegFile/_4379_ ) );
BUF_X1 \RegFile/_9230_ ( .A(\RegFile/_0266_ ), .Z(\RegFile/_4380_ ) );
BUF_X1 \RegFile/_9231_ ( .A(\RegFile/_0267_ ), .Z(\RegFile/_4381_ ) );
BUF_X1 \RegFile/_9232_ ( .A(\RegFile/_0268_ ), .Z(\RegFile/_4382_ ) );
BUF_X1 \RegFile/_9233_ ( .A(\RegFile/_0269_ ), .Z(\RegFile/_4383_ ) );
BUF_X1 \RegFile/_9234_ ( .A(\RegFile/_0270_ ), .Z(\RegFile/_4384_ ) );
BUF_X1 \RegFile/_9235_ ( .A(\RegFile/_0271_ ), .Z(\RegFile/_4385_ ) );
BUF_X1 \RegFile/_9236_ ( .A(\RegFile/_0272_ ), .Z(\RegFile/_4386_ ) );
BUF_X1 \RegFile/_9237_ ( .A(\RegFile/_0273_ ), .Z(\RegFile/_4387_ ) );
BUF_X1 \RegFile/_9238_ ( .A(\RegFile/_0274_ ), .Z(\RegFile/_4388_ ) );
BUF_X1 \RegFile/_9239_ ( .A(\RegFile/_0275_ ), .Z(\RegFile/_4389_ ) );
BUF_X1 \RegFile/_9240_ ( .A(\RegFile/_0276_ ), .Z(\RegFile/_4390_ ) );
BUF_X1 \RegFile/_9241_ ( .A(\RegFile/_0277_ ), .Z(\RegFile/_4391_ ) );
BUF_X1 \RegFile/_9242_ ( .A(\RegFile/_0278_ ), .Z(\RegFile/_4392_ ) );
BUF_X1 \RegFile/_9243_ ( .A(\RegFile/_0279_ ), .Z(\RegFile/_4393_ ) );
BUF_X1 \RegFile/_9244_ ( .A(\RegFile/_0280_ ), .Z(\RegFile/_4394_ ) );
BUF_X1 \RegFile/_9245_ ( .A(\RegFile/_0281_ ), .Z(\RegFile/_4395_ ) );
BUF_X1 \RegFile/_9246_ ( .A(\RegFile/_0282_ ), .Z(\RegFile/_4396_ ) );
BUF_X1 \RegFile/_9247_ ( .A(\RegFile/_0283_ ), .Z(\RegFile/_4397_ ) );
BUF_X1 \RegFile/_9248_ ( .A(\RegFile/_0284_ ), .Z(\RegFile/_4398_ ) );
BUF_X1 \RegFile/_9249_ ( .A(\RegFile/_0285_ ), .Z(\RegFile/_4399_ ) );
BUF_X1 \RegFile/_9250_ ( .A(\RegFile/_0286_ ), .Z(\RegFile/_4400_ ) );
BUF_X1 \RegFile/_9251_ ( .A(\RegFile/_0287_ ), .Z(\RegFile/_4401_ ) );
BUF_X1 \RegFile/_9252_ ( .A(\RegFile/_0288_ ), .Z(\RegFile/_4402_ ) );
BUF_X1 \RegFile/_9253_ ( .A(\RegFile/_0289_ ), .Z(\RegFile/_4403_ ) );
BUF_X1 \RegFile/_9254_ ( .A(\RegFile/_0290_ ), .Z(\RegFile/_4404_ ) );
BUF_X1 \RegFile/_9255_ ( .A(\RegFile/_0291_ ), .Z(\RegFile/_4405_ ) );
BUF_X1 \RegFile/_9256_ ( .A(\RegFile/_0292_ ), .Z(\RegFile/_4406_ ) );
BUF_X1 \RegFile/_9257_ ( .A(\RegFile/_0293_ ), .Z(\RegFile/_4407_ ) );
BUF_X1 \RegFile/_9258_ ( .A(\RegFile/_0294_ ), .Z(\RegFile/_4408_ ) );
BUF_X1 \RegFile/_9259_ ( .A(\RegFile/_0295_ ), .Z(\RegFile/_4409_ ) );
BUF_X1 \RegFile/_9260_ ( .A(\RegFile/_0296_ ), .Z(\RegFile/_4410_ ) );
BUF_X1 \RegFile/_9261_ ( .A(\RegFile/_0297_ ), .Z(\RegFile/_4411_ ) );
BUF_X1 \RegFile/_9262_ ( .A(\RegFile/_0298_ ), .Z(\RegFile/_4412_ ) );
BUF_X1 \RegFile/_9263_ ( .A(\RegFile/_0299_ ), .Z(\RegFile/_4413_ ) );
BUF_X1 \RegFile/_9264_ ( .A(\RegFile/_0300_ ), .Z(\RegFile/_4414_ ) );
BUF_X1 \RegFile/_9265_ ( .A(\RegFile/_0301_ ), .Z(\RegFile/_4415_ ) );
BUF_X1 \RegFile/_9266_ ( .A(\RegFile/_0302_ ), .Z(\RegFile/_4416_ ) );
BUF_X1 \RegFile/_9267_ ( .A(\RegFile/_0303_ ), .Z(\RegFile/_4417_ ) );
BUF_X1 \RegFile/_9268_ ( .A(\RegFile/_0304_ ), .Z(\RegFile/_4418_ ) );
BUF_X1 \RegFile/_9269_ ( .A(\RegFile/_0305_ ), .Z(\RegFile/_4419_ ) );
BUF_X1 \RegFile/_9270_ ( .A(\RegFile/_0306_ ), .Z(\RegFile/_4420_ ) );
BUF_X1 \RegFile/_9271_ ( .A(\RegFile/_0307_ ), .Z(\RegFile/_4421_ ) );
BUF_X1 \RegFile/_9272_ ( .A(\RegFile/_0308_ ), .Z(\RegFile/_4422_ ) );
BUF_X1 \RegFile/_9273_ ( .A(\RegFile/_0309_ ), .Z(\RegFile/_4423_ ) );
BUF_X1 \RegFile/_9274_ ( .A(\RegFile/_0310_ ), .Z(\RegFile/_4424_ ) );
BUF_X1 \RegFile/_9275_ ( .A(\RegFile/_0311_ ), .Z(\RegFile/_4425_ ) );
BUF_X1 \RegFile/_9276_ ( .A(\RegFile/_0312_ ), .Z(\RegFile/_4426_ ) );
BUF_X1 \RegFile/_9277_ ( .A(\RegFile/_0313_ ), .Z(\RegFile/_4427_ ) );
BUF_X1 \RegFile/_9278_ ( .A(\RegFile/_0314_ ), .Z(\RegFile/_4428_ ) );
BUF_X1 \RegFile/_9279_ ( .A(\RegFile/_0315_ ), .Z(\RegFile/_4429_ ) );
BUF_X1 \RegFile/_9280_ ( .A(\RegFile/_0316_ ), .Z(\RegFile/_4430_ ) );
BUF_X1 \RegFile/_9281_ ( .A(\RegFile/_0317_ ), .Z(\RegFile/_4431_ ) );
BUF_X1 \RegFile/_9282_ ( .A(\RegFile/_0318_ ), .Z(\RegFile/_4432_ ) );
BUF_X1 \RegFile/_9283_ ( .A(\RegFile/_0319_ ), .Z(\RegFile/_4433_ ) );
BUF_X1 \RegFile/_9284_ ( .A(\RegFile/_0320_ ), .Z(\RegFile/_4434_ ) );
BUF_X1 \RegFile/_9285_ ( .A(\RegFile/_0321_ ), .Z(\RegFile/_4435_ ) );
BUF_X1 \RegFile/_9286_ ( .A(\RegFile/_0322_ ), .Z(\RegFile/_4436_ ) );
BUF_X1 \RegFile/_9287_ ( .A(\RegFile/_0323_ ), .Z(\RegFile/_4437_ ) );
BUF_X1 \RegFile/_9288_ ( .A(\RegFile/_0324_ ), .Z(\RegFile/_4438_ ) );
BUF_X1 \RegFile/_9289_ ( .A(\RegFile/_0325_ ), .Z(\RegFile/_4439_ ) );
BUF_X1 \RegFile/_9290_ ( .A(\RegFile/_0326_ ), .Z(\RegFile/_4440_ ) );
BUF_X1 \RegFile/_9291_ ( .A(\RegFile/_0327_ ), .Z(\RegFile/_4441_ ) );
BUF_X1 \RegFile/_9292_ ( .A(\RegFile/_0328_ ), .Z(\RegFile/_4442_ ) );
BUF_X1 \RegFile/_9293_ ( .A(\RegFile/_0329_ ), .Z(\RegFile/_4443_ ) );
BUF_X1 \RegFile/_9294_ ( .A(\RegFile/_0330_ ), .Z(\RegFile/_4444_ ) );
BUF_X1 \RegFile/_9295_ ( .A(\RegFile/_0331_ ), .Z(\RegFile/_4445_ ) );
BUF_X1 \RegFile/_9296_ ( .A(\RegFile/_0332_ ), .Z(\RegFile/_4446_ ) );
BUF_X1 \RegFile/_9297_ ( .A(\RegFile/_0333_ ), .Z(\RegFile/_4447_ ) );
BUF_X1 \RegFile/_9298_ ( .A(\RegFile/_0334_ ), .Z(\RegFile/_4448_ ) );
BUF_X1 \RegFile/_9299_ ( .A(\RegFile/_0335_ ), .Z(\RegFile/_4449_ ) );
BUF_X1 \RegFile/_9300_ ( .A(\RegFile/_0336_ ), .Z(\RegFile/_4450_ ) );
BUF_X1 \RegFile/_9301_ ( .A(\RegFile/_0337_ ), .Z(\RegFile/_4451_ ) );
BUF_X1 \RegFile/_9302_ ( .A(\RegFile/_0338_ ), .Z(\RegFile/_4452_ ) );
BUF_X1 \RegFile/_9303_ ( .A(\RegFile/_0339_ ), .Z(\RegFile/_4453_ ) );
BUF_X1 \RegFile/_9304_ ( .A(\RegFile/_0340_ ), .Z(\RegFile/_4454_ ) );
BUF_X1 \RegFile/_9305_ ( .A(\RegFile/_0341_ ), .Z(\RegFile/_4455_ ) );
BUF_X1 \RegFile/_9306_ ( .A(\RegFile/_0342_ ), .Z(\RegFile/_4456_ ) );
BUF_X1 \RegFile/_9307_ ( .A(\RegFile/_0343_ ), .Z(\RegFile/_4457_ ) );
BUF_X1 \RegFile/_9308_ ( .A(\RegFile/_0344_ ), .Z(\RegFile/_4458_ ) );
BUF_X1 \RegFile/_9309_ ( .A(\RegFile/_0345_ ), .Z(\RegFile/_4459_ ) );
BUF_X1 \RegFile/_9310_ ( .A(\RegFile/_0346_ ), .Z(\RegFile/_4460_ ) );
BUF_X1 \RegFile/_9311_ ( .A(\RegFile/_0347_ ), .Z(\RegFile/_4461_ ) );
BUF_X1 \RegFile/_9312_ ( .A(\RegFile/_0348_ ), .Z(\RegFile/_4462_ ) );
BUF_X1 \RegFile/_9313_ ( .A(\RegFile/_0349_ ), .Z(\RegFile/_4463_ ) );
BUF_X1 \RegFile/_9314_ ( .A(\RegFile/_0350_ ), .Z(\RegFile/_4464_ ) );
BUF_X1 \RegFile/_9315_ ( .A(\RegFile/_0351_ ), .Z(\RegFile/_4465_ ) );
BUF_X1 \RegFile/_9316_ ( .A(\RegFile/_0352_ ), .Z(\RegFile/_4466_ ) );
BUF_X1 \RegFile/_9317_ ( .A(\RegFile/_0353_ ), .Z(\RegFile/_4467_ ) );
BUF_X1 \RegFile/_9318_ ( .A(\RegFile/_0354_ ), .Z(\RegFile/_4468_ ) );
BUF_X1 \RegFile/_9319_ ( .A(\RegFile/_0355_ ), .Z(\RegFile/_4469_ ) );
BUF_X1 \RegFile/_9320_ ( .A(\RegFile/_0356_ ), .Z(\RegFile/_4470_ ) );
BUF_X1 \RegFile/_9321_ ( .A(\RegFile/_0357_ ), .Z(\RegFile/_4471_ ) );
BUF_X1 \RegFile/_9322_ ( .A(\RegFile/_0358_ ), .Z(\RegFile/_4472_ ) );
BUF_X1 \RegFile/_9323_ ( .A(\RegFile/_0359_ ), .Z(\RegFile/_4473_ ) );
BUF_X1 \RegFile/_9324_ ( .A(\RegFile/_0360_ ), .Z(\RegFile/_4474_ ) );
BUF_X1 \RegFile/_9325_ ( .A(\RegFile/_0361_ ), .Z(\RegFile/_4475_ ) );
BUF_X1 \RegFile/_9326_ ( .A(\RegFile/_0362_ ), .Z(\RegFile/_4476_ ) );
BUF_X1 \RegFile/_9327_ ( .A(\RegFile/_0363_ ), .Z(\RegFile/_4477_ ) );
BUF_X1 \RegFile/_9328_ ( .A(\RegFile/_0364_ ), .Z(\RegFile/_4478_ ) );
BUF_X1 \RegFile/_9329_ ( .A(\RegFile/_0365_ ), .Z(\RegFile/_4479_ ) );
BUF_X1 \RegFile/_9330_ ( .A(\RegFile/_0366_ ), .Z(\RegFile/_4480_ ) );
BUF_X1 \RegFile/_9331_ ( .A(\RegFile/_0367_ ), .Z(\RegFile/_4481_ ) );
BUF_X1 \RegFile/_9332_ ( .A(\RegFile/_0368_ ), .Z(\RegFile/_4482_ ) );
BUF_X1 \RegFile/_9333_ ( .A(\RegFile/_0369_ ), .Z(\RegFile/_4483_ ) );
BUF_X1 \RegFile/_9334_ ( .A(\RegFile/_0370_ ), .Z(\RegFile/_4484_ ) );
BUF_X1 \RegFile/_9335_ ( .A(\RegFile/_0371_ ), .Z(\RegFile/_4485_ ) );
BUF_X1 \RegFile/_9336_ ( .A(\RegFile/_0372_ ), .Z(\RegFile/_4486_ ) );
BUF_X1 \RegFile/_9337_ ( .A(\RegFile/_0373_ ), .Z(\RegFile/_4487_ ) );
BUF_X1 \RegFile/_9338_ ( .A(\RegFile/_0374_ ), .Z(\RegFile/_4488_ ) );
BUF_X1 \RegFile/_9339_ ( .A(\RegFile/_0375_ ), .Z(\RegFile/_4489_ ) );
BUF_X1 \RegFile/_9340_ ( .A(\RegFile/_0376_ ), .Z(\RegFile/_4490_ ) );
BUF_X1 \RegFile/_9341_ ( .A(\RegFile/_0377_ ), .Z(\RegFile/_4491_ ) );
BUF_X1 \RegFile/_9342_ ( .A(\RegFile/_0378_ ), .Z(\RegFile/_4492_ ) );
BUF_X1 \RegFile/_9343_ ( .A(\RegFile/_0379_ ), .Z(\RegFile/_4493_ ) );
BUF_X1 \RegFile/_9344_ ( .A(\RegFile/_0380_ ), .Z(\RegFile/_4494_ ) );
BUF_X1 \RegFile/_9345_ ( .A(\RegFile/_0381_ ), .Z(\RegFile/_4495_ ) );
BUF_X1 \RegFile/_9346_ ( .A(\RegFile/_0382_ ), .Z(\RegFile/_4496_ ) );
BUF_X1 \RegFile/_9347_ ( .A(\RegFile/_0383_ ), .Z(\RegFile/_4497_ ) );
BUF_X1 \RegFile/_9348_ ( .A(\RegFile/_0384_ ), .Z(\RegFile/_4498_ ) );
BUF_X1 \RegFile/_9349_ ( .A(\RegFile/_0385_ ), .Z(\RegFile/_4499_ ) );
BUF_X1 \RegFile/_9350_ ( .A(\RegFile/_0386_ ), .Z(\RegFile/_4500_ ) );
BUF_X1 \RegFile/_9351_ ( .A(\RegFile/_0387_ ), .Z(\RegFile/_4501_ ) );
BUF_X1 \RegFile/_9352_ ( .A(\RegFile/_0388_ ), .Z(\RegFile/_4502_ ) );
BUF_X1 \RegFile/_9353_ ( .A(\RegFile/_0389_ ), .Z(\RegFile/_4503_ ) );
BUF_X1 \RegFile/_9354_ ( .A(\RegFile/_0390_ ), .Z(\RegFile/_4504_ ) );
BUF_X1 \RegFile/_9355_ ( .A(\RegFile/_0391_ ), .Z(\RegFile/_4505_ ) );
BUF_X1 \RegFile/_9356_ ( .A(\RegFile/_0392_ ), .Z(\RegFile/_4506_ ) );
BUF_X1 \RegFile/_9357_ ( .A(\RegFile/_0393_ ), .Z(\RegFile/_4507_ ) );
BUF_X1 \RegFile/_9358_ ( .A(\RegFile/_0394_ ), .Z(\RegFile/_4508_ ) );
BUF_X1 \RegFile/_9359_ ( .A(\RegFile/_0395_ ), .Z(\RegFile/_4509_ ) );
BUF_X1 \RegFile/_9360_ ( .A(\RegFile/_0396_ ), .Z(\RegFile/_4510_ ) );
BUF_X1 \RegFile/_9361_ ( .A(\RegFile/_0397_ ), .Z(\RegFile/_4511_ ) );
BUF_X1 \RegFile/_9362_ ( .A(\RegFile/_0398_ ), .Z(\RegFile/_4512_ ) );
BUF_X1 \RegFile/_9363_ ( .A(\RegFile/_0399_ ), .Z(\RegFile/_4513_ ) );
BUF_X1 \RegFile/_9364_ ( .A(\RegFile/_0400_ ), .Z(\RegFile/_4514_ ) );
BUF_X1 \RegFile/_9365_ ( .A(\RegFile/_0401_ ), .Z(\RegFile/_4515_ ) );
BUF_X1 \RegFile/_9366_ ( .A(\RegFile/_0402_ ), .Z(\RegFile/_4516_ ) );
BUF_X1 \RegFile/_9367_ ( .A(\RegFile/_0403_ ), .Z(\RegFile/_4517_ ) );
BUF_X1 \RegFile/_9368_ ( .A(\RegFile/_0404_ ), .Z(\RegFile/_4518_ ) );
BUF_X1 \RegFile/_9369_ ( .A(\RegFile/_0405_ ), .Z(\RegFile/_4519_ ) );
BUF_X1 \RegFile/_9370_ ( .A(\RegFile/_0406_ ), .Z(\RegFile/_4520_ ) );
BUF_X1 \RegFile/_9371_ ( .A(\RegFile/_0407_ ), .Z(\RegFile/_4521_ ) );
BUF_X1 \RegFile/_9372_ ( .A(\RegFile/_0408_ ), .Z(\RegFile/_4522_ ) );
BUF_X1 \RegFile/_9373_ ( .A(\RegFile/_0409_ ), .Z(\RegFile/_4523_ ) );
BUF_X1 \RegFile/_9374_ ( .A(\RegFile/_0410_ ), .Z(\RegFile/_4524_ ) );
BUF_X1 \RegFile/_9375_ ( .A(\RegFile/_0411_ ), .Z(\RegFile/_4525_ ) );
BUF_X1 \RegFile/_9376_ ( .A(\RegFile/_0412_ ), .Z(\RegFile/_4526_ ) );
BUF_X1 \RegFile/_9377_ ( .A(\RegFile/_0413_ ), .Z(\RegFile/_4527_ ) );
BUF_X1 \RegFile/_9378_ ( .A(\RegFile/_0414_ ), .Z(\RegFile/_4528_ ) );
BUF_X1 \RegFile/_9379_ ( .A(\RegFile/_0415_ ), .Z(\RegFile/_4529_ ) );
BUF_X1 \RegFile/_9380_ ( .A(\RegFile/_0416_ ), .Z(\RegFile/_4530_ ) );
BUF_X1 \RegFile/_9381_ ( .A(\RegFile/_0417_ ), .Z(\RegFile/_4531_ ) );
BUF_X1 \RegFile/_9382_ ( .A(\RegFile/_0418_ ), .Z(\RegFile/_4532_ ) );
BUF_X1 \RegFile/_9383_ ( .A(\RegFile/_0419_ ), .Z(\RegFile/_4533_ ) );
BUF_X1 \RegFile/_9384_ ( .A(\RegFile/_0420_ ), .Z(\RegFile/_4534_ ) );
BUF_X1 \RegFile/_9385_ ( .A(\RegFile/_0421_ ), .Z(\RegFile/_4535_ ) );
BUF_X1 \RegFile/_9386_ ( .A(\RegFile/_0422_ ), .Z(\RegFile/_4536_ ) );
BUF_X1 \RegFile/_9387_ ( .A(\RegFile/_0423_ ), .Z(\RegFile/_4537_ ) );
BUF_X1 \RegFile/_9388_ ( .A(\RegFile/_0424_ ), .Z(\RegFile/_4538_ ) );
BUF_X1 \RegFile/_9389_ ( .A(\RegFile/_0425_ ), .Z(\RegFile/_4539_ ) );
BUF_X1 \RegFile/_9390_ ( .A(\RegFile/_0426_ ), .Z(\RegFile/_4540_ ) );
BUF_X1 \RegFile/_9391_ ( .A(\RegFile/_0427_ ), .Z(\RegFile/_4541_ ) );
BUF_X1 \RegFile/_9392_ ( .A(\RegFile/_0428_ ), .Z(\RegFile/_4542_ ) );
BUF_X1 \RegFile/_9393_ ( .A(\RegFile/_0429_ ), .Z(\RegFile/_4543_ ) );
BUF_X1 \RegFile/_9394_ ( .A(\RegFile/_0430_ ), .Z(\RegFile/_4544_ ) );
BUF_X1 \RegFile/_9395_ ( .A(\RegFile/_0431_ ), .Z(\RegFile/_4545_ ) );
BUF_X1 \RegFile/_9396_ ( .A(\RegFile/_0432_ ), .Z(\RegFile/_4546_ ) );
BUF_X1 \RegFile/_9397_ ( .A(\RegFile/_0433_ ), .Z(\RegFile/_4547_ ) );
BUF_X1 \RegFile/_9398_ ( .A(\RegFile/_0434_ ), .Z(\RegFile/_4548_ ) );
BUF_X1 \RegFile/_9399_ ( .A(\RegFile/_0435_ ), .Z(\RegFile/_4549_ ) );
BUF_X1 \RegFile/_9400_ ( .A(\RegFile/_0436_ ), .Z(\RegFile/_4550_ ) );
BUF_X1 \RegFile/_9401_ ( .A(\RegFile/_0437_ ), .Z(\RegFile/_4551_ ) );
BUF_X1 \RegFile/_9402_ ( .A(\RegFile/_0438_ ), .Z(\RegFile/_4552_ ) );
BUF_X1 \RegFile/_9403_ ( .A(\RegFile/_0439_ ), .Z(\RegFile/_4553_ ) );
BUF_X1 \RegFile/_9404_ ( .A(\RegFile/_0440_ ), .Z(\RegFile/_4554_ ) );
BUF_X1 \RegFile/_9405_ ( .A(\RegFile/_0441_ ), .Z(\RegFile/_4555_ ) );
BUF_X1 \RegFile/_9406_ ( .A(\RegFile/_0442_ ), .Z(\RegFile/_4556_ ) );
BUF_X1 \RegFile/_9407_ ( .A(\RegFile/_0443_ ), .Z(\RegFile/_4557_ ) );
BUF_X1 \RegFile/_9408_ ( .A(\RegFile/_0444_ ), .Z(\RegFile/_4558_ ) );
BUF_X1 \RegFile/_9409_ ( .A(\RegFile/_0445_ ), .Z(\RegFile/_4559_ ) );
BUF_X1 \RegFile/_9410_ ( .A(\RegFile/_0446_ ), .Z(\RegFile/_4560_ ) );
BUF_X1 \RegFile/_9411_ ( .A(\RegFile/_0447_ ), .Z(\RegFile/_4561_ ) );
BUF_X1 \RegFile/_9412_ ( .A(\RegFile/_0448_ ), .Z(\RegFile/_4562_ ) );
BUF_X1 \RegFile/_9413_ ( .A(\RegFile/_0449_ ), .Z(\RegFile/_4563_ ) );
BUF_X1 \RegFile/_9414_ ( .A(\RegFile/_0450_ ), .Z(\RegFile/_4564_ ) );
BUF_X1 \RegFile/_9415_ ( .A(\RegFile/_0451_ ), .Z(\RegFile/_4565_ ) );
BUF_X1 \RegFile/_9416_ ( .A(\RegFile/_0452_ ), .Z(\RegFile/_4566_ ) );
BUF_X1 \RegFile/_9417_ ( .A(\RegFile/_0453_ ), .Z(\RegFile/_4567_ ) );
BUF_X1 \RegFile/_9418_ ( .A(\RegFile/_0454_ ), .Z(\RegFile/_4568_ ) );
BUF_X1 \RegFile/_9419_ ( .A(\RegFile/_0455_ ), .Z(\RegFile/_4569_ ) );
BUF_X1 \RegFile/_9420_ ( .A(\RegFile/_0456_ ), .Z(\RegFile/_4570_ ) );
BUF_X1 \RegFile/_9421_ ( .A(\RegFile/_0457_ ), .Z(\RegFile/_4571_ ) );
BUF_X1 \RegFile/_9422_ ( .A(\RegFile/_0458_ ), .Z(\RegFile/_4572_ ) );
BUF_X1 \RegFile/_9423_ ( .A(\RegFile/_0459_ ), .Z(\RegFile/_4573_ ) );
BUF_X1 \RegFile/_9424_ ( .A(\RegFile/_0460_ ), .Z(\RegFile/_4574_ ) );
BUF_X1 \RegFile/_9425_ ( .A(\RegFile/_0461_ ), .Z(\RegFile/_4575_ ) );
BUF_X1 \RegFile/_9426_ ( .A(\RegFile/_0462_ ), .Z(\RegFile/_4576_ ) );
BUF_X1 \RegFile/_9427_ ( .A(\RegFile/_0463_ ), .Z(\RegFile/_4577_ ) );
BUF_X1 \RegFile/_9428_ ( .A(\RegFile/_0464_ ), .Z(\RegFile/_4578_ ) );
BUF_X1 \RegFile/_9429_ ( .A(\RegFile/_0465_ ), .Z(\RegFile/_4579_ ) );
BUF_X1 \RegFile/_9430_ ( .A(\RegFile/_0466_ ), .Z(\RegFile/_4580_ ) );
BUF_X1 \RegFile/_9431_ ( .A(\RegFile/_0467_ ), .Z(\RegFile/_4581_ ) );
BUF_X1 \RegFile/_9432_ ( .A(\RegFile/_0468_ ), .Z(\RegFile/_4582_ ) );
BUF_X1 \RegFile/_9433_ ( .A(\RegFile/_0469_ ), .Z(\RegFile/_4583_ ) );
BUF_X1 \RegFile/_9434_ ( .A(\RegFile/_0470_ ), .Z(\RegFile/_4584_ ) );
BUF_X1 \RegFile/_9435_ ( .A(\RegFile/_0471_ ), .Z(\RegFile/_4585_ ) );
BUF_X1 \RegFile/_9436_ ( .A(\RegFile/_0472_ ), .Z(\RegFile/_4586_ ) );
BUF_X1 \RegFile/_9437_ ( .A(\RegFile/_0473_ ), .Z(\RegFile/_4587_ ) );
BUF_X1 \RegFile/_9438_ ( .A(\RegFile/_0474_ ), .Z(\RegFile/_4588_ ) );
BUF_X1 \RegFile/_9439_ ( .A(\RegFile/_0475_ ), .Z(\RegFile/_4589_ ) );
BUF_X1 \RegFile/_9440_ ( .A(\RegFile/_0476_ ), .Z(\RegFile/_4590_ ) );
BUF_X1 \RegFile/_9441_ ( .A(\RegFile/_0477_ ), .Z(\RegFile/_4591_ ) );
BUF_X1 \RegFile/_9442_ ( .A(\RegFile/_0478_ ), .Z(\RegFile/_4592_ ) );
BUF_X1 \RegFile/_9443_ ( .A(\RegFile/_0479_ ), .Z(\RegFile/_4593_ ) );
BUF_X1 \RegFile/_9444_ ( .A(\RegFile/_0480_ ), .Z(\RegFile/_4594_ ) );
BUF_X1 \RegFile/_9445_ ( .A(\RegFile/_0481_ ), .Z(\RegFile/_4595_ ) );
BUF_X1 \RegFile/_9446_ ( .A(\RegFile/_0482_ ), .Z(\RegFile/_4596_ ) );
BUF_X1 \RegFile/_9447_ ( .A(\RegFile/_0483_ ), .Z(\RegFile/_4597_ ) );
BUF_X1 \RegFile/_9448_ ( .A(\RegFile/_0484_ ), .Z(\RegFile/_4598_ ) );
BUF_X1 \RegFile/_9449_ ( .A(\RegFile/_0485_ ), .Z(\RegFile/_4599_ ) );
BUF_X1 \RegFile/_9450_ ( .A(\RegFile/_0486_ ), .Z(\RegFile/_4600_ ) );
BUF_X1 \RegFile/_9451_ ( .A(\RegFile/_0487_ ), .Z(\RegFile/_4601_ ) );
BUF_X1 \RegFile/_9452_ ( .A(\RegFile/_0488_ ), .Z(\RegFile/_4602_ ) );
BUF_X1 \RegFile/_9453_ ( .A(\RegFile/_0489_ ), .Z(\RegFile/_4603_ ) );
BUF_X1 \RegFile/_9454_ ( .A(\RegFile/_0490_ ), .Z(\RegFile/_4604_ ) );
BUF_X1 \RegFile/_9455_ ( .A(\RegFile/_0491_ ), .Z(\RegFile/_4605_ ) );
BUF_X1 \RegFile/_9456_ ( .A(\RegFile/_0492_ ), .Z(\RegFile/_4606_ ) );
BUF_X1 \RegFile/_9457_ ( .A(\RegFile/_0493_ ), .Z(\RegFile/_4607_ ) );
BUF_X1 \RegFile/_9458_ ( .A(\RegFile/_0494_ ), .Z(\RegFile/_4608_ ) );
BUF_X1 \RegFile/_9459_ ( .A(\RegFile/_0495_ ), .Z(\RegFile/_4609_ ) );
BUF_X1 \RegFile/_9460_ ( .A(\RegFile/_0496_ ), .Z(\RegFile/_4610_ ) );
BUF_X1 \RegFile/_9461_ ( .A(\RegFile/_0497_ ), .Z(\RegFile/_4611_ ) );
BUF_X1 \RegFile/_9462_ ( .A(\RegFile/_0498_ ), .Z(\RegFile/_4612_ ) );
BUF_X1 \RegFile/_9463_ ( .A(\RegFile/_0499_ ), .Z(\RegFile/_4613_ ) );
BUF_X1 \RegFile/_9464_ ( .A(\RegFile/_0500_ ), .Z(\RegFile/_4614_ ) );
BUF_X1 \RegFile/_9465_ ( .A(\RegFile/_0501_ ), .Z(\RegFile/_4615_ ) );
BUF_X1 \RegFile/_9466_ ( .A(\RegFile/_0502_ ), .Z(\RegFile/_4616_ ) );
BUF_X1 \RegFile/_9467_ ( .A(\RegFile/_0503_ ), .Z(\RegFile/_4617_ ) );
BUF_X1 \RegFile/_9468_ ( .A(\RegFile/_0504_ ), .Z(\RegFile/_4618_ ) );
BUF_X1 \RegFile/_9469_ ( .A(\RegFile/_0505_ ), .Z(\RegFile/_4619_ ) );
BUF_X1 \RegFile/_9470_ ( .A(\RegFile/_0506_ ), .Z(\RegFile/_4620_ ) );
BUF_X1 \RegFile/_9471_ ( .A(\RegFile/_0507_ ), .Z(\RegFile/_4621_ ) );
BUF_X1 \RegFile/_9472_ ( .A(\RegFile/_0508_ ), .Z(\RegFile/_4622_ ) );
BUF_X1 \RegFile/_9473_ ( .A(\RegFile/_0509_ ), .Z(\RegFile/_4623_ ) );
BUF_X1 \RegFile/_9474_ ( .A(\RegFile/_0510_ ), .Z(\RegFile/_4624_ ) );
BUF_X1 \RegFile/_9475_ ( .A(\RegFile/_0511_ ), .Z(\RegFile/_4625_ ) );
BUF_X1 \RegFile/_9476_ ( .A(\RegFile/_0512_ ), .Z(\RegFile/_4626_ ) );
BUF_X1 \RegFile/_9477_ ( .A(\RegFile/_0513_ ), .Z(\RegFile/_4627_ ) );
BUF_X1 \RegFile/_9478_ ( .A(\RegFile/_0514_ ), .Z(\RegFile/_4628_ ) );
BUF_X1 \RegFile/_9479_ ( .A(\RegFile/_0515_ ), .Z(\RegFile/_4629_ ) );
BUF_X1 \RegFile/_9480_ ( .A(\RegFile/_0516_ ), .Z(\RegFile/_4630_ ) );
BUF_X1 \RegFile/_9481_ ( .A(\RegFile/_0517_ ), .Z(\RegFile/_4631_ ) );
BUF_X1 \RegFile/_9482_ ( .A(\RegFile/_0518_ ), .Z(\RegFile/_4632_ ) );
BUF_X1 \RegFile/_9483_ ( .A(\RegFile/_0519_ ), .Z(\RegFile/_4633_ ) );
BUF_X1 \RegFile/_9484_ ( .A(\RegFile/_0520_ ), .Z(\RegFile/_4634_ ) );
BUF_X1 \RegFile/_9485_ ( .A(\RegFile/_0521_ ), .Z(\RegFile/_4635_ ) );
BUF_X1 \RegFile/_9486_ ( .A(\RegFile/_0522_ ), .Z(\RegFile/_4636_ ) );
BUF_X1 \RegFile/_9487_ ( .A(\RegFile/_0523_ ), .Z(\RegFile/_4637_ ) );
BUF_X1 \RegFile/_9488_ ( .A(\RegFile/_0524_ ), .Z(\RegFile/_4638_ ) );
BUF_X1 \RegFile/_9489_ ( .A(\RegFile/_0525_ ), .Z(\RegFile/_4639_ ) );
BUF_X1 \RegFile/_9490_ ( .A(\RegFile/_0526_ ), .Z(\RegFile/_4640_ ) );
BUF_X1 \RegFile/_9491_ ( .A(\RegFile/_0527_ ), .Z(\RegFile/_4641_ ) );
BUF_X1 \RegFile/_9492_ ( .A(\RegFile/_0528_ ), .Z(\RegFile/_4642_ ) );
BUF_X1 \RegFile/_9493_ ( .A(\RegFile/_0529_ ), .Z(\RegFile/_4643_ ) );
BUF_X1 \RegFile/_9494_ ( .A(\RegFile/_0530_ ), .Z(\RegFile/_4644_ ) );
BUF_X1 \RegFile/_9495_ ( .A(\RegFile/_0531_ ), .Z(\RegFile/_4645_ ) );
BUF_X1 \RegFile/_9496_ ( .A(\RegFile/_0532_ ), .Z(\RegFile/_4646_ ) );
BUF_X1 \RegFile/_9497_ ( .A(\RegFile/_0533_ ), .Z(\RegFile/_4647_ ) );
BUF_X1 \RegFile/_9498_ ( .A(\RegFile/_0534_ ), .Z(\RegFile/_4648_ ) );
BUF_X1 \RegFile/_9499_ ( .A(\RegFile/_0535_ ), .Z(\RegFile/_4649_ ) );
BUF_X1 \RegFile/_9500_ ( .A(\RegFile/_0536_ ), .Z(\RegFile/_4650_ ) );
BUF_X1 \RegFile/_9501_ ( .A(\RegFile/_0537_ ), .Z(\RegFile/_4651_ ) );
BUF_X1 \RegFile/_9502_ ( .A(\RegFile/_0538_ ), .Z(\RegFile/_4652_ ) );
BUF_X1 \RegFile/_9503_ ( .A(\RegFile/_0539_ ), .Z(\RegFile/_4653_ ) );
BUF_X1 \RegFile/_9504_ ( .A(\RegFile/_0540_ ), .Z(\RegFile/_4654_ ) );
BUF_X1 \RegFile/_9505_ ( .A(\RegFile/_0541_ ), .Z(\RegFile/_4655_ ) );
BUF_X1 \RegFile/_9506_ ( .A(\RegFile/_0542_ ), .Z(\RegFile/_4656_ ) );
BUF_X1 \RegFile/_9507_ ( .A(\RegFile/_0543_ ), .Z(\RegFile/_4657_ ) );
BUF_X1 \RegFile/_9508_ ( .A(\RegFile/_0544_ ), .Z(\RegFile/_4658_ ) );
BUF_X1 \RegFile/_9509_ ( .A(\RegFile/_0545_ ), .Z(\RegFile/_4659_ ) );
BUF_X1 \RegFile/_9510_ ( .A(\RegFile/_0546_ ), .Z(\RegFile/_4660_ ) );
BUF_X1 \RegFile/_9511_ ( .A(\RegFile/_0547_ ), .Z(\RegFile/_4661_ ) );
BUF_X1 \RegFile/_9512_ ( .A(\RegFile/_0548_ ), .Z(\RegFile/_4662_ ) );
BUF_X1 \RegFile/_9513_ ( .A(\RegFile/_0549_ ), .Z(\RegFile/_4663_ ) );
BUF_X1 \RegFile/_9514_ ( .A(\RegFile/_0550_ ), .Z(\RegFile/_4664_ ) );
BUF_X1 \RegFile/_9515_ ( .A(\RegFile/_0551_ ), .Z(\RegFile/_4665_ ) );
BUF_X1 \RegFile/_9516_ ( .A(\RegFile/_0552_ ), .Z(\RegFile/_4666_ ) );
BUF_X1 \RegFile/_9517_ ( .A(\RegFile/_0553_ ), .Z(\RegFile/_4667_ ) );
BUF_X1 \RegFile/_9518_ ( .A(\RegFile/_0554_ ), .Z(\RegFile/_4668_ ) );
BUF_X1 \RegFile/_9519_ ( .A(\RegFile/_0555_ ), .Z(\RegFile/_4669_ ) );
BUF_X1 \RegFile/_9520_ ( .A(\RegFile/_0556_ ), .Z(\RegFile/_4670_ ) );
BUF_X1 \RegFile/_9521_ ( .A(\RegFile/_0557_ ), .Z(\RegFile/_4671_ ) );
BUF_X1 \RegFile/_9522_ ( .A(\RegFile/_0558_ ), .Z(\RegFile/_4672_ ) );
BUF_X1 \RegFile/_9523_ ( .A(\RegFile/_0559_ ), .Z(\RegFile/_4673_ ) );
BUF_X1 \RegFile/_9524_ ( .A(\RegFile/_0560_ ), .Z(\RegFile/_4674_ ) );
BUF_X1 \RegFile/_9525_ ( .A(\RegFile/_0561_ ), .Z(\RegFile/_4675_ ) );
BUF_X1 \RegFile/_9526_ ( .A(\RegFile/_0562_ ), .Z(\RegFile/_4676_ ) );
BUF_X1 \RegFile/_9527_ ( .A(\RegFile/_0563_ ), .Z(\RegFile/_4677_ ) );
BUF_X1 \RegFile/_9528_ ( .A(\RegFile/_0564_ ), .Z(\RegFile/_4678_ ) );
BUF_X1 \RegFile/_9529_ ( .A(\RegFile/_0565_ ), .Z(\RegFile/_4679_ ) );
BUF_X1 \RegFile/_9530_ ( .A(\RegFile/_0566_ ), .Z(\RegFile/_4680_ ) );
BUF_X1 \RegFile/_9531_ ( .A(\RegFile/_0567_ ), .Z(\RegFile/_4681_ ) );
BUF_X1 \RegFile/_9532_ ( .A(\RegFile/_0568_ ), .Z(\RegFile/_4682_ ) );
BUF_X1 \RegFile/_9533_ ( .A(\RegFile/_0569_ ), .Z(\RegFile/_4683_ ) );
BUF_X1 \RegFile/_9534_ ( .A(\RegFile/_0570_ ), .Z(\RegFile/_4684_ ) );
BUF_X1 \RegFile/_9535_ ( .A(\RegFile/_0571_ ), .Z(\RegFile/_4685_ ) );
BUF_X1 \RegFile/_9536_ ( .A(\RegFile/_0572_ ), .Z(\RegFile/_4686_ ) );
BUF_X1 \RegFile/_9537_ ( .A(\RegFile/_0573_ ), .Z(\RegFile/_4687_ ) );
BUF_X1 \RegFile/_9538_ ( .A(\RegFile/_0574_ ), .Z(\RegFile/_4688_ ) );
BUF_X1 \RegFile/_9539_ ( .A(\RegFile/_0575_ ), .Z(\RegFile/_4689_ ) );
BUF_X1 \RegFile/_9540_ ( .A(\RegFile/_0576_ ), .Z(\RegFile/_4690_ ) );
BUF_X1 \RegFile/_9541_ ( .A(\RegFile/_0577_ ), .Z(\RegFile/_4691_ ) );
BUF_X1 \RegFile/_9542_ ( .A(\RegFile/_0578_ ), .Z(\RegFile/_4692_ ) );
BUF_X1 \RegFile/_9543_ ( .A(\RegFile/_0579_ ), .Z(\RegFile/_4693_ ) );
BUF_X1 \RegFile/_9544_ ( .A(\RegFile/_0580_ ), .Z(\RegFile/_4694_ ) );
BUF_X1 \RegFile/_9545_ ( .A(\RegFile/_0581_ ), .Z(\RegFile/_4695_ ) );
BUF_X1 \RegFile/_9546_ ( .A(\RegFile/_0582_ ), .Z(\RegFile/_4696_ ) );
BUF_X1 \RegFile/_9547_ ( .A(\RegFile/_0583_ ), .Z(\RegFile/_4697_ ) );
BUF_X1 \RegFile/_9548_ ( .A(\RegFile/_0584_ ), .Z(\RegFile/_4698_ ) );
BUF_X1 \RegFile/_9549_ ( .A(\RegFile/_0585_ ), .Z(\RegFile/_4699_ ) );
BUF_X1 \RegFile/_9550_ ( .A(\RegFile/_0586_ ), .Z(\RegFile/_4700_ ) );
BUF_X1 \RegFile/_9551_ ( .A(\RegFile/_0587_ ), .Z(\RegFile/_4701_ ) );
BUF_X1 \RegFile/_9552_ ( .A(\RegFile/_0588_ ), .Z(\RegFile/_4702_ ) );
BUF_X1 \RegFile/_9553_ ( .A(\RegFile/_0589_ ), .Z(\RegFile/_4703_ ) );
BUF_X1 \RegFile/_9554_ ( .A(\RegFile/_0590_ ), .Z(\RegFile/_4704_ ) );
BUF_X1 \RegFile/_9555_ ( .A(\RegFile/_0591_ ), .Z(\RegFile/_4705_ ) );
BUF_X1 \RegFile/_9556_ ( .A(\RegFile/_0592_ ), .Z(\RegFile/_4706_ ) );
BUF_X1 \RegFile/_9557_ ( .A(\RegFile/_0593_ ), .Z(\RegFile/_4707_ ) );
BUF_X1 \RegFile/_9558_ ( .A(\RegFile/_0594_ ), .Z(\RegFile/_4708_ ) );
BUF_X1 \RegFile/_9559_ ( .A(\RegFile/_0595_ ), .Z(\RegFile/_4709_ ) );
BUF_X1 \RegFile/_9560_ ( .A(\RegFile/_0596_ ), .Z(\RegFile/_4710_ ) );
BUF_X1 \RegFile/_9561_ ( .A(\RegFile/_0597_ ), .Z(\RegFile/_4711_ ) );
BUF_X1 \RegFile/_9562_ ( .A(\RegFile/_0598_ ), .Z(\RegFile/_4712_ ) );
BUF_X1 \RegFile/_9563_ ( .A(\RegFile/_0599_ ), .Z(\RegFile/_4713_ ) );
BUF_X1 \RegFile/_9564_ ( .A(\RegFile/_0600_ ), .Z(\RegFile/_4714_ ) );
BUF_X1 \RegFile/_9565_ ( .A(\RegFile/_0601_ ), .Z(\RegFile/_4715_ ) );
BUF_X1 \RegFile/_9566_ ( .A(\RegFile/_0602_ ), .Z(\RegFile/_4716_ ) );
BUF_X1 \RegFile/_9567_ ( .A(\RegFile/_0603_ ), .Z(\RegFile/_4717_ ) );
BUF_X1 \RegFile/_9568_ ( .A(\RegFile/_0604_ ), .Z(\RegFile/_4718_ ) );
BUF_X1 \RegFile/_9569_ ( .A(\RegFile/_0605_ ), .Z(\RegFile/_4719_ ) );
BUF_X1 \RegFile/_9570_ ( .A(\RegFile/_0606_ ), .Z(\RegFile/_4720_ ) );
BUF_X1 \RegFile/_9571_ ( .A(\RegFile/_0607_ ), .Z(\RegFile/_4721_ ) );
MUX2_X1 \WBU/_275_ ( .A(\WBU/_133_ ), .B(\WBU/_069_ ), .S(fanout_net_20 ), .Z(\WBU/_166_ ) );
MUX2_X1 \WBU/_276_ ( .A(\WBU/_144_ ), .B(\WBU/_080_ ), .S(fanout_net_20 ), .Z(\WBU/_177_ ) );
MUX2_X1 \WBU/_277_ ( .A(\WBU/_155_ ), .B(\WBU/_091_ ), .S(fanout_net_20 ), .Z(\WBU/_188_ ) );
MUX2_X1 \WBU/_278_ ( .A(\WBU/_158_ ), .B(\WBU/_094_ ), .S(fanout_net_20 ), .Z(\WBU/_191_ ) );
MUX2_X1 \WBU/_279_ ( .A(\WBU/_159_ ), .B(\WBU/_095_ ), .S(fanout_net_20 ), .Z(\WBU/_192_ ) );
MUX2_X1 \WBU/_280_ ( .A(\WBU/_160_ ), .B(\WBU/_096_ ), .S(fanout_net_20 ), .Z(\WBU/_193_ ) );
MUX2_X1 \WBU/_281_ ( .A(\WBU/_161_ ), .B(\WBU/_097_ ), .S(fanout_net_20 ), .Z(\WBU/_194_ ) );
MUX2_X1 \WBU/_282_ ( .A(\WBU/_162_ ), .B(\WBU/_098_ ), .S(fanout_net_20 ), .Z(\WBU/_195_ ) );
MUX2_X1 \WBU/_283_ ( .A(\WBU/_163_ ), .B(\WBU/_099_ ), .S(fanout_net_20 ), .Z(\WBU/_196_ ) );
MUX2_X1 \WBU/_284_ ( .A(\WBU/_164_ ), .B(\WBU/_100_ ), .S(fanout_net_20 ), .Z(\WBU/_197_ ) );
MUX2_X1 \WBU/_285_ ( .A(\WBU/_134_ ), .B(\WBU/_070_ ), .S(fanout_net_20 ), .Z(\WBU/_167_ ) );
MUX2_X1 \WBU/_286_ ( .A(\WBU/_135_ ), .B(\WBU/_071_ ), .S(fanout_net_20 ), .Z(\WBU/_168_ ) );
MUX2_X1 \WBU/_287_ ( .A(\WBU/_136_ ), .B(\WBU/_072_ ), .S(fanout_net_20 ), .Z(\WBU/_169_ ) );
MUX2_X1 \WBU/_288_ ( .A(\WBU/_137_ ), .B(\WBU/_073_ ), .S(fanout_net_20 ), .Z(\WBU/_170_ ) );
MUX2_X1 \WBU/_289_ ( .A(\WBU/_138_ ), .B(\WBU/_074_ ), .S(fanout_net_20 ), .Z(\WBU/_171_ ) );
MUX2_X1 \WBU/_290_ ( .A(\WBU/_139_ ), .B(\WBU/_075_ ), .S(fanout_net_20 ), .Z(\WBU/_172_ ) );
MUX2_X1 \WBU/_291_ ( .A(\WBU/_140_ ), .B(\WBU/_076_ ), .S(fanout_net_20 ), .Z(\WBU/_173_ ) );
MUX2_X1 \WBU/_292_ ( .A(\WBU/_141_ ), .B(\WBU/_077_ ), .S(fanout_net_20 ), .Z(\WBU/_174_ ) );
MUX2_X1 \WBU/_293_ ( .A(\WBU/_142_ ), .B(\WBU/_078_ ), .S(fanout_net_20 ), .Z(\WBU/_175_ ) );
MUX2_X1 \WBU/_294_ ( .A(\WBU/_143_ ), .B(\WBU/_079_ ), .S(fanout_net_20 ), .Z(\WBU/_176_ ) );
MUX2_X1 \WBU/_295_ ( .A(\WBU/_145_ ), .B(\WBU/_081_ ), .S(fanout_net_20 ), .Z(\WBU/_178_ ) );
MUX2_X1 \WBU/_296_ ( .A(\WBU/_146_ ), .B(\WBU/_082_ ), .S(fanout_net_20 ), .Z(\WBU/_179_ ) );
MUX2_X1 \WBU/_297_ ( .A(\WBU/_147_ ), .B(\WBU/_083_ ), .S(fanout_net_20 ), .Z(\WBU/_180_ ) );
MUX2_X1 \WBU/_298_ ( .A(\WBU/_148_ ), .B(\WBU/_084_ ), .S(fanout_net_20 ), .Z(\WBU/_181_ ) );
MUX2_X1 \WBU/_299_ ( .A(\WBU/_149_ ), .B(\WBU/_085_ ), .S(fanout_net_20 ), .Z(\WBU/_182_ ) );
MUX2_X1 \WBU/_300_ ( .A(\WBU/_150_ ), .B(\WBU/_086_ ), .S(fanout_net_20 ), .Z(\WBU/_183_ ) );
MUX2_X1 \WBU/_301_ ( .A(\WBU/_151_ ), .B(\WBU/_087_ ), .S(fanout_net_20 ), .Z(\WBU/_184_ ) );
MUX2_X1 \WBU/_302_ ( .A(\WBU/_152_ ), .B(\WBU/_088_ ), .S(fanout_net_20 ), .Z(\WBU/_185_ ) );
MUX2_X1 \WBU/_303_ ( .A(\WBU/_153_ ), .B(\WBU/_089_ ), .S(fanout_net_20 ), .Z(\WBU/_186_ ) );
MUX2_X1 \WBU/_304_ ( .A(\WBU/_154_ ), .B(\WBU/_090_ ), .S(fanout_net_20 ), .Z(\WBU/_187_ ) );
MUX2_X1 \WBU/_305_ ( .A(\WBU/_156_ ), .B(\WBU/_092_ ), .S(\WBU/_065_ ), .Z(\WBU/_189_ ) );
MUX2_X1 \WBU/_306_ ( .A(\WBU/_157_ ), .B(\WBU/_093_ ), .S(\WBU/_065_ ), .Z(\WBU/_190_ ) );
INV_X32 \WBU/_307_ ( .A(\WBU/_067_ ), .ZN(\WBU/_198_ ) );
AND2_X2 \WBU/_308_ ( .A1(\WBU/_198_ ), .A2(\WBU/_068_ ), .ZN(\WBU/_199_ ) );
BUF_X8 \WBU/_309_ ( .A(\WBU/_199_ ), .Z(\WBU/_200_ ) );
NOR2_X4 \WBU/_310_ ( .A1(\WBU/_198_ ), .A2(\WBU/_068_ ), .ZN(\WBU/_201_ ) );
BUF_X4 \WBU/_311_ ( .A(\WBU/_201_ ), .Z(\WBU/_202_ ) );
AOI22_X1 \WBU/_312_ ( .A1(\WBU/_200_ ), .A2(\WBU/_069_ ), .B1(\WBU/_202_ ), .B2(\WBU/_101_ ), .ZN(\WBU/_203_ ) );
XNOR2_X2 \WBU/_313_ ( .A(\WBU/_067_ ), .B(\WBU/_068_ ), .ZN(\WBU/_204_ ) );
BUF_X4 \WBU/_314_ ( .A(\WBU/_204_ ), .Z(\WBU/_205_ ) );
NAND2_X1 \WBU/_315_ ( .A1(\WBU/_205_ ), .A2(\WBU/_033_ ), .ZN(\WBU/_206_ ) );
NAND2_X1 \WBU/_316_ ( .A1(\WBU/_203_ ), .A2(\WBU/_206_ ), .ZN(\WBU/_000_ ) );
AOI22_X1 \WBU/_317_ ( .A1(\WBU/_200_ ), .A2(\WBU/_080_ ), .B1(\WBU/_202_ ), .B2(\WBU/_112_ ), .ZN(\WBU/_207_ ) );
NAND2_X1 \WBU/_318_ ( .A1(\WBU/_205_ ), .A2(\WBU/_044_ ), .ZN(\WBU/_208_ ) );
NAND2_X1 \WBU/_319_ ( .A1(\WBU/_207_ ), .A2(\WBU/_208_ ), .ZN(\WBU/_011_ ) );
AOI22_X1 \WBU/_320_ ( .A1(\WBU/_200_ ), .A2(\WBU/_091_ ), .B1(\WBU/_202_ ), .B2(\WBU/_123_ ), .ZN(\WBU/_209_ ) );
NAND2_X1 \WBU/_321_ ( .A1(\WBU/_205_ ), .A2(\WBU/_055_ ), .ZN(\WBU/_210_ ) );
NAND2_X1 \WBU/_322_ ( .A1(\WBU/_209_ ), .A2(\WBU/_210_ ), .ZN(\WBU/_022_ ) );
AOI22_X1 \WBU/_323_ ( .A1(\WBU/_200_ ), .A2(\WBU/_094_ ), .B1(\WBU/_202_ ), .B2(\WBU/_126_ ), .ZN(\WBU/_211_ ) );
NAND2_X1 \WBU/_324_ ( .A1(\WBU/_205_ ), .A2(\WBU/_058_ ), .ZN(\WBU/_212_ ) );
NAND2_X1 \WBU/_325_ ( .A1(\WBU/_211_ ), .A2(\WBU/_212_ ), .ZN(\WBU/_025_ ) );
AOI22_X1 \WBU/_326_ ( .A1(\WBU/_200_ ), .A2(\WBU/_095_ ), .B1(\WBU/_202_ ), .B2(\WBU/_127_ ), .ZN(\WBU/_213_ ) );
NAND2_X1 \WBU/_327_ ( .A1(\WBU/_205_ ), .A2(\WBU/_059_ ), .ZN(\WBU/_214_ ) );
NAND2_X1 \WBU/_328_ ( .A1(\WBU/_213_ ), .A2(\WBU/_214_ ), .ZN(\WBU/_026_ ) );
AOI22_X1 \WBU/_329_ ( .A1(\WBU/_200_ ), .A2(\WBU/_096_ ), .B1(\WBU/_202_ ), .B2(\WBU/_128_ ), .ZN(\WBU/_215_ ) );
NAND2_X1 \WBU/_330_ ( .A1(\WBU/_205_ ), .A2(\WBU/_060_ ), .ZN(\WBU/_216_ ) );
NAND2_X1 \WBU/_331_ ( .A1(\WBU/_215_ ), .A2(\WBU/_216_ ), .ZN(\WBU/_027_ ) );
AOI22_X1 \WBU/_332_ ( .A1(\WBU/_200_ ), .A2(\WBU/_097_ ), .B1(\WBU/_202_ ), .B2(\WBU/_129_ ), .ZN(\WBU/_217_ ) );
NAND2_X1 \WBU/_333_ ( .A1(\WBU/_205_ ), .A2(\WBU/_061_ ), .ZN(\WBU/_218_ ) );
NAND2_X1 \WBU/_334_ ( .A1(\WBU/_217_ ), .A2(\WBU/_218_ ), .ZN(\WBU/_028_ ) );
AOI22_X1 \WBU/_335_ ( .A1(\WBU/_200_ ), .A2(\WBU/_098_ ), .B1(\WBU/_202_ ), .B2(\WBU/_130_ ), .ZN(\WBU/_219_ ) );
NAND2_X1 \WBU/_336_ ( .A1(\WBU/_205_ ), .A2(\WBU/_062_ ), .ZN(\WBU/_220_ ) );
NAND2_X1 \WBU/_337_ ( .A1(\WBU/_219_ ), .A2(\WBU/_220_ ), .ZN(\WBU/_029_ ) );
AOI22_X1 \WBU/_338_ ( .A1(\WBU/_200_ ), .A2(\WBU/_099_ ), .B1(\WBU/_202_ ), .B2(\WBU/_131_ ), .ZN(\WBU/_221_ ) );
NAND2_X1 \WBU/_339_ ( .A1(\WBU/_205_ ), .A2(\WBU/_063_ ), .ZN(\WBU/_222_ ) );
NAND2_X1 \WBU/_340_ ( .A1(\WBU/_221_ ), .A2(\WBU/_222_ ), .ZN(\WBU/_030_ ) );
AOI22_X1 \WBU/_341_ ( .A1(\WBU/_200_ ), .A2(\WBU/_100_ ), .B1(\WBU/_202_ ), .B2(\WBU/_132_ ), .ZN(\WBU/_223_ ) );
NAND2_X1 \WBU/_342_ ( .A1(\WBU/_205_ ), .A2(\WBU/_064_ ), .ZN(\WBU/_224_ ) );
NAND2_X1 \WBU/_343_ ( .A1(\WBU/_223_ ), .A2(\WBU/_224_ ), .ZN(\WBU/_031_ ) );
BUF_X8 \WBU/_344_ ( .A(\WBU/_199_ ), .Z(\WBU/_225_ ) );
BUF_X4 \WBU/_345_ ( .A(\WBU/_201_ ), .Z(\WBU/_226_ ) );
AOI22_X1 \WBU/_346_ ( .A1(\WBU/_225_ ), .A2(\WBU/_070_ ), .B1(\WBU/_226_ ), .B2(\WBU/_102_ ), .ZN(\WBU/_227_ ) );
BUF_X4 \WBU/_347_ ( .A(\WBU/_204_ ), .Z(\WBU/_228_ ) );
NAND2_X1 \WBU/_348_ ( .A1(\WBU/_228_ ), .A2(\WBU/_034_ ), .ZN(\WBU/_229_ ) );
NAND2_X1 \WBU/_349_ ( .A1(\WBU/_227_ ), .A2(\WBU/_229_ ), .ZN(\WBU/_001_ ) );
AOI22_X1 \WBU/_350_ ( .A1(\WBU/_225_ ), .A2(\WBU/_071_ ), .B1(\WBU/_226_ ), .B2(\WBU/_103_ ), .ZN(\WBU/_230_ ) );
NAND2_X1 \WBU/_351_ ( .A1(\WBU/_228_ ), .A2(\WBU/_035_ ), .ZN(\WBU/_231_ ) );
NAND2_X1 \WBU/_352_ ( .A1(\WBU/_230_ ), .A2(\WBU/_231_ ), .ZN(\WBU/_002_ ) );
AOI22_X1 \WBU/_353_ ( .A1(\WBU/_225_ ), .A2(\WBU/_072_ ), .B1(\WBU/_226_ ), .B2(\WBU/_104_ ), .ZN(\WBU/_232_ ) );
NAND2_X1 \WBU/_354_ ( .A1(\WBU/_228_ ), .A2(\WBU/_036_ ), .ZN(\WBU/_233_ ) );
NAND2_X1 \WBU/_355_ ( .A1(\WBU/_232_ ), .A2(\WBU/_233_ ), .ZN(\WBU/_003_ ) );
AOI22_X1 \WBU/_356_ ( .A1(\WBU/_225_ ), .A2(\WBU/_073_ ), .B1(\WBU/_226_ ), .B2(\WBU/_105_ ), .ZN(\WBU/_234_ ) );
NAND2_X1 \WBU/_357_ ( .A1(\WBU/_228_ ), .A2(\WBU/_037_ ), .ZN(\WBU/_235_ ) );
NAND2_X1 \WBU/_358_ ( .A1(\WBU/_234_ ), .A2(\WBU/_235_ ), .ZN(\WBU/_004_ ) );
AOI22_X1 \WBU/_359_ ( .A1(\WBU/_225_ ), .A2(\WBU/_074_ ), .B1(\WBU/_226_ ), .B2(\WBU/_106_ ), .ZN(\WBU/_236_ ) );
NAND2_X1 \WBU/_360_ ( .A1(\WBU/_228_ ), .A2(\WBU/_038_ ), .ZN(\WBU/_237_ ) );
NAND2_X1 \WBU/_361_ ( .A1(\WBU/_236_ ), .A2(\WBU/_237_ ), .ZN(\WBU/_005_ ) );
AOI22_X1 \WBU/_362_ ( .A1(\WBU/_225_ ), .A2(\WBU/_075_ ), .B1(\WBU/_226_ ), .B2(\WBU/_107_ ), .ZN(\WBU/_238_ ) );
NAND2_X1 \WBU/_363_ ( .A1(\WBU/_228_ ), .A2(\WBU/_039_ ), .ZN(\WBU/_239_ ) );
NAND2_X1 \WBU/_364_ ( .A1(\WBU/_238_ ), .A2(\WBU/_239_ ), .ZN(\WBU/_006_ ) );
AOI22_X1 \WBU/_365_ ( .A1(\WBU/_225_ ), .A2(\WBU/_076_ ), .B1(\WBU/_226_ ), .B2(\WBU/_108_ ), .ZN(\WBU/_240_ ) );
NAND2_X1 \WBU/_366_ ( .A1(\WBU/_228_ ), .A2(\WBU/_040_ ), .ZN(\WBU/_241_ ) );
NAND2_X1 \WBU/_367_ ( .A1(\WBU/_240_ ), .A2(\WBU/_241_ ), .ZN(\WBU/_007_ ) );
AOI22_X1 \WBU/_368_ ( .A1(\WBU/_225_ ), .A2(\WBU/_077_ ), .B1(\WBU/_226_ ), .B2(\WBU/_109_ ), .ZN(\WBU/_242_ ) );
NAND2_X1 \WBU/_369_ ( .A1(\WBU/_228_ ), .A2(\WBU/_041_ ), .ZN(\WBU/_243_ ) );
NAND2_X1 \WBU/_370_ ( .A1(\WBU/_242_ ), .A2(\WBU/_243_ ), .ZN(\WBU/_008_ ) );
AOI22_X1 \WBU/_371_ ( .A1(\WBU/_225_ ), .A2(\WBU/_078_ ), .B1(\WBU/_226_ ), .B2(\WBU/_110_ ), .ZN(\WBU/_244_ ) );
NAND2_X1 \WBU/_372_ ( .A1(\WBU/_228_ ), .A2(\WBU/_042_ ), .ZN(\WBU/_245_ ) );
NAND2_X1 \WBU/_373_ ( .A1(\WBU/_244_ ), .A2(\WBU/_245_ ), .ZN(\WBU/_009_ ) );
AOI22_X1 \WBU/_374_ ( .A1(\WBU/_225_ ), .A2(\WBU/_079_ ), .B1(\WBU/_226_ ), .B2(\WBU/_111_ ), .ZN(\WBU/_246_ ) );
NAND2_X1 \WBU/_375_ ( .A1(\WBU/_228_ ), .A2(\WBU/_043_ ), .ZN(\WBU/_247_ ) );
NAND2_X1 \WBU/_376_ ( .A1(\WBU/_246_ ), .A2(\WBU/_247_ ), .ZN(\WBU/_010_ ) );
BUF_X8 \WBU/_377_ ( .A(\WBU/_199_ ), .Z(\WBU/_248_ ) );
BUF_X4 \WBU/_378_ ( .A(\WBU/_201_ ), .Z(\WBU/_249_ ) );
AOI22_X1 \WBU/_379_ ( .A1(\WBU/_248_ ), .A2(\WBU/_081_ ), .B1(\WBU/_249_ ), .B2(\WBU/_113_ ), .ZN(\WBU/_250_ ) );
BUF_X4 \WBU/_380_ ( .A(\WBU/_204_ ), .Z(\WBU/_251_ ) );
NAND2_X1 \WBU/_381_ ( .A1(\WBU/_251_ ), .A2(\WBU/_045_ ), .ZN(\WBU/_252_ ) );
NAND2_X1 \WBU/_382_ ( .A1(\WBU/_250_ ), .A2(\WBU/_252_ ), .ZN(\WBU/_012_ ) );
AOI22_X1 \WBU/_383_ ( .A1(\WBU/_248_ ), .A2(\WBU/_082_ ), .B1(\WBU/_249_ ), .B2(\WBU/_114_ ), .ZN(\WBU/_253_ ) );
NAND2_X1 \WBU/_384_ ( .A1(\WBU/_251_ ), .A2(\WBU/_046_ ), .ZN(\WBU/_254_ ) );
NAND2_X1 \WBU/_385_ ( .A1(\WBU/_253_ ), .A2(\WBU/_254_ ), .ZN(\WBU/_013_ ) );
AOI22_X1 \WBU/_386_ ( .A1(\WBU/_248_ ), .A2(\WBU/_083_ ), .B1(\WBU/_249_ ), .B2(\WBU/_115_ ), .ZN(\WBU/_255_ ) );
NAND2_X1 \WBU/_387_ ( .A1(\WBU/_251_ ), .A2(\WBU/_047_ ), .ZN(\WBU/_256_ ) );
NAND2_X1 \WBU/_388_ ( .A1(\WBU/_255_ ), .A2(\WBU/_256_ ), .ZN(\WBU/_014_ ) );
AOI22_X1 \WBU/_389_ ( .A1(\WBU/_248_ ), .A2(\WBU/_084_ ), .B1(\WBU/_249_ ), .B2(\WBU/_116_ ), .ZN(\WBU/_257_ ) );
NAND2_X1 \WBU/_390_ ( .A1(\WBU/_251_ ), .A2(\WBU/_048_ ), .ZN(\WBU/_258_ ) );
NAND2_X1 \WBU/_391_ ( .A1(\WBU/_257_ ), .A2(\WBU/_258_ ), .ZN(\WBU/_015_ ) );
AOI22_X1 \WBU/_392_ ( .A1(\WBU/_248_ ), .A2(\WBU/_085_ ), .B1(\WBU/_249_ ), .B2(\WBU/_117_ ), .ZN(\WBU/_259_ ) );
NAND2_X1 \WBU/_393_ ( .A1(\WBU/_251_ ), .A2(\WBU/_049_ ), .ZN(\WBU/_260_ ) );
NAND2_X1 \WBU/_394_ ( .A1(\WBU/_259_ ), .A2(\WBU/_260_ ), .ZN(\WBU/_016_ ) );
AOI22_X1 \WBU/_395_ ( .A1(\WBU/_248_ ), .A2(\WBU/_086_ ), .B1(\WBU/_249_ ), .B2(\WBU/_118_ ), .ZN(\WBU/_261_ ) );
NAND2_X1 \WBU/_396_ ( .A1(\WBU/_251_ ), .A2(\WBU/_050_ ), .ZN(\WBU/_262_ ) );
NAND2_X1 \WBU/_397_ ( .A1(\WBU/_261_ ), .A2(\WBU/_262_ ), .ZN(\WBU/_017_ ) );
AOI22_X1 \WBU/_398_ ( .A1(\WBU/_248_ ), .A2(\WBU/_087_ ), .B1(\WBU/_249_ ), .B2(\WBU/_119_ ), .ZN(\WBU/_263_ ) );
NAND2_X1 \WBU/_399_ ( .A1(\WBU/_251_ ), .A2(\WBU/_051_ ), .ZN(\WBU/_264_ ) );
NAND2_X1 \WBU/_400_ ( .A1(\WBU/_263_ ), .A2(\WBU/_264_ ), .ZN(\WBU/_018_ ) );
AOI22_X1 \WBU/_401_ ( .A1(\WBU/_248_ ), .A2(\WBU/_088_ ), .B1(\WBU/_249_ ), .B2(\WBU/_120_ ), .ZN(\WBU/_265_ ) );
NAND2_X1 \WBU/_402_ ( .A1(\WBU/_251_ ), .A2(\WBU/_052_ ), .ZN(\WBU/_266_ ) );
NAND2_X1 \WBU/_403_ ( .A1(\WBU/_265_ ), .A2(\WBU/_266_ ), .ZN(\WBU/_019_ ) );
AOI22_X1 \WBU/_404_ ( .A1(\WBU/_248_ ), .A2(\WBU/_089_ ), .B1(\WBU/_249_ ), .B2(\WBU/_121_ ), .ZN(\WBU/_267_ ) );
NAND2_X1 \WBU/_405_ ( .A1(\WBU/_251_ ), .A2(\WBU/_053_ ), .ZN(\WBU/_268_ ) );
NAND2_X1 \WBU/_406_ ( .A1(\WBU/_267_ ), .A2(\WBU/_268_ ), .ZN(\WBU/_020_ ) );
AOI22_X1 \WBU/_407_ ( .A1(\WBU/_248_ ), .A2(\WBU/_090_ ), .B1(\WBU/_249_ ), .B2(\WBU/_122_ ), .ZN(\WBU/_269_ ) );
NAND2_X1 \WBU/_408_ ( .A1(\WBU/_251_ ), .A2(\WBU/_054_ ), .ZN(\WBU/_270_ ) );
NAND2_X1 \WBU/_409_ ( .A1(\WBU/_269_ ), .A2(\WBU/_270_ ), .ZN(\WBU/_021_ ) );
AOI22_X1 \WBU/_410_ ( .A1(\WBU/_199_ ), .A2(\WBU/_092_ ), .B1(\WBU/_201_ ), .B2(\WBU/_124_ ), .ZN(\WBU/_271_ ) );
NAND2_X1 \WBU/_411_ ( .A1(\WBU/_204_ ), .A2(\WBU/_056_ ), .ZN(\WBU/_272_ ) );
NAND2_X1 \WBU/_412_ ( .A1(\WBU/_271_ ), .A2(\WBU/_272_ ), .ZN(\WBU/_023_ ) );
AOI22_X1 \WBU/_413_ ( .A1(\WBU/_199_ ), .A2(\WBU/_093_ ), .B1(\WBU/_201_ ), .B2(\WBU/_125_ ), .ZN(\WBU/_273_ ) );
NAND2_X1 \WBU/_414_ ( .A1(\WBU/_204_ ), .A2(\WBU/_057_ ), .ZN(\WBU/_274_ ) );
NAND2_X1 \WBU/_415_ ( .A1(\WBU/_273_ ), .A2(\WBU/_274_ ), .ZN(\WBU/_024_ ) );
AND2_X1 \WBU/_416_ ( .A1(\WBU/_165_ ), .A2(\WBU/_066_ ), .ZN(\WBU/_032_ ) );
BUF_X1 \WBU/_417_ ( .A(\_EXU_io_out_bits_wa [0] ), .Z(\_WBU_io_RegFileAccess_wa [0] ) );
BUF_X1 \WBU/_418_ ( .A(\_EXU_io_out_bits_wa [1] ), .Z(\_WBU_io_RegFileAccess_wa [1] ) );
BUF_X1 \WBU/_419_ ( .A(\_EXU_io_out_bits_wa [2] ), .Z(\_WBU_io_RegFileAccess_wa [2] ) );
BUF_X1 \WBU/_420_ ( .A(\_EXU_io_out_bits_wa [3] ), .Z(\_WBU_io_RegFileAccess_wa [3] ) );
BUF_X1 \WBU/_421_ ( .A(_IFU_io_in_ready ), .Z(_WBU_io_in_ready ) );
BUF_X1 \WBU/_422_ ( .A(_EXU_io_out_valid ), .Z(_WBU_io_out_valid ) );
BUF_X1 \WBU/_423_ ( .A(\_EXU_io_out_bits_pcCom [0] ), .Z(\WBU/_133_ ) );
BUF_X1 \WBU/_424_ ( .A(\_EXU_io_out_bits_csrOut [0] ), .Z(\WBU/_069_ ) );
BUF_X1 \WBU/_425_ ( .A(_EXU_io_out_bits_control_pcSrc ), .Z(\WBU/_065_ ) );
BUF_X1 \WBU/_426_ ( .A(\WBU/_166_ ), .Z(\_WBU_io_out_bits_nextPc [0] ) );
BUF_X1 \WBU/_427_ ( .A(\_EXU_io_out_bits_pcCom [1] ), .Z(\WBU/_144_ ) );
BUF_X1 \WBU/_428_ ( .A(\_EXU_io_out_bits_csrOut [1] ), .Z(\WBU/_080_ ) );
BUF_X1 \WBU/_429_ ( .A(\WBU/_177_ ), .Z(\_WBU_io_out_bits_nextPc [1] ) );
BUF_X1 \WBU/_430_ ( .A(\_EXU_io_out_bits_pcCom [2] ), .Z(\WBU/_155_ ) );
BUF_X1 \WBU/_431_ ( .A(\_EXU_io_out_bits_csrOut [2] ), .Z(\WBU/_091_ ) );
BUF_X1 \WBU/_432_ ( .A(\WBU/_188_ ), .Z(\_WBU_io_out_bits_nextPc [2] ) );
BUF_X1 \WBU/_433_ ( .A(\_EXU_io_out_bits_pcCom [3] ), .Z(\WBU/_158_ ) );
BUF_X1 \WBU/_434_ ( .A(\_EXU_io_out_bits_csrOut [3] ), .Z(\WBU/_094_ ) );
BUF_X1 \WBU/_435_ ( .A(\WBU/_191_ ), .Z(\_WBU_io_out_bits_nextPc [3] ) );
BUF_X1 \WBU/_436_ ( .A(\_EXU_io_out_bits_pcCom [4] ), .Z(\WBU/_159_ ) );
BUF_X1 \WBU/_437_ ( .A(\_EXU_io_out_bits_csrOut [4] ), .Z(\WBU/_095_ ) );
BUF_X1 \WBU/_438_ ( .A(\WBU/_192_ ), .Z(\_WBU_io_out_bits_nextPc [4] ) );
BUF_X1 \WBU/_439_ ( .A(\_EXU_io_out_bits_pcCom [5] ), .Z(\WBU/_160_ ) );
BUF_X1 \WBU/_440_ ( .A(\_EXU_io_out_bits_csrOut [5] ), .Z(\WBU/_096_ ) );
BUF_X1 \WBU/_441_ ( .A(\WBU/_193_ ), .Z(\_WBU_io_out_bits_nextPc [5] ) );
BUF_X1 \WBU/_442_ ( .A(\_EXU_io_out_bits_pcCom [6] ), .Z(\WBU/_161_ ) );
BUF_X1 \WBU/_443_ ( .A(\_EXU_io_out_bits_csrOut [6] ), .Z(\WBU/_097_ ) );
BUF_X1 \WBU/_444_ ( .A(\WBU/_194_ ), .Z(\_WBU_io_out_bits_nextPc [6] ) );
BUF_X1 \WBU/_445_ ( .A(\_EXU_io_out_bits_pcCom [7] ), .Z(\WBU/_162_ ) );
BUF_X1 \WBU/_446_ ( .A(\_EXU_io_out_bits_csrOut [7] ), .Z(\WBU/_098_ ) );
BUF_X1 \WBU/_447_ ( .A(\WBU/_195_ ), .Z(\_WBU_io_out_bits_nextPc [7] ) );
BUF_X1 \WBU/_448_ ( .A(\_EXU_io_out_bits_pcCom [8] ), .Z(\WBU/_163_ ) );
BUF_X1 \WBU/_449_ ( .A(\_EXU_io_out_bits_csrOut [8] ), .Z(\WBU/_099_ ) );
BUF_X1 \WBU/_450_ ( .A(\WBU/_196_ ), .Z(\_WBU_io_out_bits_nextPc [8] ) );
BUF_X1 \WBU/_451_ ( .A(\_EXU_io_out_bits_pcCom [9] ), .Z(\WBU/_164_ ) );
BUF_X1 \WBU/_452_ ( .A(\_EXU_io_out_bits_csrOut [9] ), .Z(\WBU/_100_ ) );
BUF_X1 \WBU/_453_ ( .A(\WBU/_197_ ), .Z(\_WBU_io_out_bits_nextPc [9] ) );
BUF_X1 \WBU/_454_ ( .A(\_EXU_io_out_bits_pcCom [10] ), .Z(\WBU/_134_ ) );
BUF_X1 \WBU/_455_ ( .A(\_EXU_io_out_bits_csrOut [10] ), .Z(\WBU/_070_ ) );
BUF_X1 \WBU/_456_ ( .A(\WBU/_167_ ), .Z(\_WBU_io_out_bits_nextPc [10] ) );
BUF_X1 \WBU/_457_ ( .A(\_EXU_io_out_bits_pcCom [11] ), .Z(\WBU/_135_ ) );
BUF_X1 \WBU/_458_ ( .A(\_EXU_io_out_bits_csrOut [11] ), .Z(\WBU/_071_ ) );
BUF_X1 \WBU/_459_ ( .A(\WBU/_168_ ), .Z(\_WBU_io_out_bits_nextPc [11] ) );
BUF_X1 \WBU/_460_ ( .A(\_EXU_io_out_bits_pcCom [12] ), .Z(\WBU/_136_ ) );
BUF_X1 \WBU/_461_ ( .A(\_EXU_io_out_bits_csrOut [12] ), .Z(\WBU/_072_ ) );
BUF_X1 \WBU/_462_ ( .A(\WBU/_169_ ), .Z(\_WBU_io_out_bits_nextPc [12] ) );
BUF_X1 \WBU/_463_ ( .A(\_EXU_io_out_bits_pcCom [13] ), .Z(\WBU/_137_ ) );
BUF_X1 \WBU/_464_ ( .A(\_EXU_io_out_bits_csrOut [13] ), .Z(\WBU/_073_ ) );
BUF_X1 \WBU/_465_ ( .A(\WBU/_170_ ), .Z(\_WBU_io_out_bits_nextPc [13] ) );
BUF_X1 \WBU/_466_ ( .A(\_EXU_io_out_bits_pcCom [14] ), .Z(\WBU/_138_ ) );
BUF_X1 \WBU/_467_ ( .A(\_EXU_io_out_bits_csrOut [14] ), .Z(\WBU/_074_ ) );
BUF_X1 \WBU/_468_ ( .A(\WBU/_171_ ), .Z(\_WBU_io_out_bits_nextPc [14] ) );
BUF_X1 \WBU/_469_ ( .A(\_EXU_io_out_bits_pcCom [15] ), .Z(\WBU/_139_ ) );
BUF_X1 \WBU/_470_ ( .A(\_EXU_io_out_bits_csrOut [15] ), .Z(\WBU/_075_ ) );
BUF_X1 \WBU/_471_ ( .A(\WBU/_172_ ), .Z(\_WBU_io_out_bits_nextPc [15] ) );
BUF_X1 \WBU/_472_ ( .A(\_EXU_io_out_bits_pcCom [16] ), .Z(\WBU/_140_ ) );
BUF_X1 \WBU/_473_ ( .A(\_EXU_io_out_bits_csrOut [16] ), .Z(\WBU/_076_ ) );
BUF_X1 \WBU/_474_ ( .A(\WBU/_173_ ), .Z(\_WBU_io_out_bits_nextPc [16] ) );
BUF_X1 \WBU/_475_ ( .A(\_EXU_io_out_bits_pcCom [17] ), .Z(\WBU/_141_ ) );
BUF_X1 \WBU/_476_ ( .A(\_EXU_io_out_bits_csrOut [17] ), .Z(\WBU/_077_ ) );
BUF_X1 \WBU/_477_ ( .A(\WBU/_174_ ), .Z(\_WBU_io_out_bits_nextPc [17] ) );
BUF_X1 \WBU/_478_ ( .A(\_EXU_io_out_bits_pcCom [18] ), .Z(\WBU/_142_ ) );
BUF_X1 \WBU/_479_ ( .A(\_EXU_io_out_bits_csrOut [18] ), .Z(\WBU/_078_ ) );
BUF_X1 \WBU/_480_ ( .A(\WBU/_175_ ), .Z(\_WBU_io_out_bits_nextPc [18] ) );
BUF_X1 \WBU/_481_ ( .A(\_EXU_io_out_bits_pcCom [19] ), .Z(\WBU/_143_ ) );
BUF_X1 \WBU/_482_ ( .A(\_EXU_io_out_bits_csrOut [19] ), .Z(\WBU/_079_ ) );
BUF_X1 \WBU/_483_ ( .A(\WBU/_176_ ), .Z(\_WBU_io_out_bits_nextPc [19] ) );
BUF_X1 \WBU/_484_ ( .A(\_EXU_io_out_bits_pcCom [20] ), .Z(\WBU/_145_ ) );
BUF_X1 \WBU/_485_ ( .A(\_EXU_io_out_bits_csrOut [20] ), .Z(\WBU/_081_ ) );
BUF_X1 \WBU/_486_ ( .A(\WBU/_178_ ), .Z(\_WBU_io_out_bits_nextPc [20] ) );
BUF_X1 \WBU/_487_ ( .A(\_EXU_io_out_bits_pcCom [21] ), .Z(\WBU/_146_ ) );
BUF_X1 \WBU/_488_ ( .A(\_EXU_io_out_bits_csrOut [21] ), .Z(\WBU/_082_ ) );
BUF_X1 \WBU/_489_ ( .A(\WBU/_179_ ), .Z(\_WBU_io_out_bits_nextPc [21] ) );
BUF_X1 \WBU/_490_ ( .A(\_EXU_io_out_bits_pcCom [22] ), .Z(\WBU/_147_ ) );
BUF_X1 \WBU/_491_ ( .A(\_EXU_io_out_bits_csrOut [22] ), .Z(\WBU/_083_ ) );
BUF_X1 \WBU/_492_ ( .A(\WBU/_180_ ), .Z(\_WBU_io_out_bits_nextPc [22] ) );
BUF_X1 \WBU/_493_ ( .A(\_EXU_io_out_bits_pcCom [23] ), .Z(\WBU/_148_ ) );
BUF_X1 \WBU/_494_ ( .A(\_EXU_io_out_bits_csrOut [23] ), .Z(\WBU/_084_ ) );
BUF_X1 \WBU/_495_ ( .A(\WBU/_181_ ), .Z(\_WBU_io_out_bits_nextPc [23] ) );
BUF_X1 \WBU/_496_ ( .A(\_EXU_io_out_bits_pcCom [24] ), .Z(\WBU/_149_ ) );
BUF_X1 \WBU/_497_ ( .A(\_EXU_io_out_bits_csrOut [24] ), .Z(\WBU/_085_ ) );
BUF_X1 \WBU/_498_ ( .A(\WBU/_182_ ), .Z(\_WBU_io_out_bits_nextPc [24] ) );
BUF_X1 \WBU/_499_ ( .A(\_EXU_io_out_bits_pcCom [25] ), .Z(\WBU/_150_ ) );
BUF_X1 \WBU/_500_ ( .A(\_EXU_io_out_bits_csrOut [25] ), .Z(\WBU/_086_ ) );
BUF_X1 \WBU/_501_ ( .A(\WBU/_183_ ), .Z(\_WBU_io_out_bits_nextPc [25] ) );
BUF_X1 \WBU/_502_ ( .A(\_EXU_io_out_bits_pcCom [26] ), .Z(\WBU/_151_ ) );
BUF_X1 \WBU/_503_ ( .A(\_EXU_io_out_bits_csrOut [26] ), .Z(\WBU/_087_ ) );
BUF_X1 \WBU/_504_ ( .A(\WBU/_184_ ), .Z(\_WBU_io_out_bits_nextPc [26] ) );
BUF_X1 \WBU/_505_ ( .A(\_EXU_io_out_bits_pcCom [27] ), .Z(\WBU/_152_ ) );
BUF_X1 \WBU/_506_ ( .A(\_EXU_io_out_bits_csrOut [27] ), .Z(\WBU/_088_ ) );
BUF_X1 \WBU/_507_ ( .A(\WBU/_185_ ), .Z(\_WBU_io_out_bits_nextPc [27] ) );
BUF_X1 \WBU/_508_ ( .A(\_EXU_io_out_bits_pcCom [28] ), .Z(\WBU/_153_ ) );
BUF_X1 \WBU/_509_ ( .A(\_EXU_io_out_bits_csrOut [28] ), .Z(\WBU/_089_ ) );
BUF_X1 \WBU/_510_ ( .A(\WBU/_186_ ), .Z(\_WBU_io_out_bits_nextPc [28] ) );
BUF_X1 \WBU/_511_ ( .A(\_EXU_io_out_bits_pcCom [29] ), .Z(\WBU/_154_ ) );
BUF_X1 \WBU/_512_ ( .A(\_EXU_io_out_bits_csrOut [29] ), .Z(\WBU/_090_ ) );
BUF_X1 \WBU/_513_ ( .A(\WBU/_187_ ), .Z(\_WBU_io_out_bits_nextPc [29] ) );
BUF_X1 \WBU/_514_ ( .A(\_EXU_io_out_bits_pcCom [30] ), .Z(\WBU/_156_ ) );
BUF_X1 \WBU/_515_ ( .A(\_EXU_io_out_bits_csrOut [30] ), .Z(\WBU/_092_ ) );
BUF_X1 \WBU/_516_ ( .A(\WBU/_189_ ), .Z(\_WBU_io_out_bits_nextPc [30] ) );
BUF_X1 \WBU/_517_ ( .A(\_EXU_io_out_bits_pcCom [31] ), .Z(\WBU/_157_ ) );
BUF_X1 \WBU/_518_ ( .A(\_EXU_io_out_bits_csrOut [31] ), .Z(\WBU/_093_ ) );
BUF_X1 \WBU/_519_ ( .A(\WBU/_190_ ), .Z(\_WBU_io_out_bits_nextPc [31] ) );
BUF_X1 \WBU/_520_ ( .A(\_EXU_io_out_bits_control_wbSrc [0] ), .Z(\WBU/_067_ ) );
BUF_X1 \WBU/_521_ ( .A(\_EXU_io_out_bits_control_wbSrc [1] ), .Z(\WBU/_068_ ) );
BUF_X1 \WBU/_522_ ( .A(\_EXU_io_out_bits_memOut [0] ), .Z(\WBU/_101_ ) );
BUF_X1 \WBU/_523_ ( .A(\_EXU_io_out_bits_aluOut [0] ), .Z(\WBU/_033_ ) );
BUF_X1 \WBU/_524_ ( .A(\WBU/_000_ ), .Z(\_WBU_io_RegFileAccess_wd [0] ) );
BUF_X1 \WBU/_525_ ( .A(\_EXU_io_out_bits_memOut [1] ), .Z(\WBU/_112_ ) );
BUF_X1 \WBU/_526_ ( .A(\_EXU_io_out_bits_aluOut [1] ), .Z(\WBU/_044_ ) );
BUF_X1 \WBU/_527_ ( .A(\WBU/_011_ ), .Z(\_WBU_io_RegFileAccess_wd [1] ) );
BUF_X1 \WBU/_528_ ( .A(\_EXU_io_out_bits_memOut [2] ), .Z(\WBU/_123_ ) );
BUF_X1 \WBU/_529_ ( .A(\_EXU_io_out_bits_aluOut [2] ), .Z(\WBU/_055_ ) );
BUF_X1 \WBU/_530_ ( .A(\WBU/_022_ ), .Z(\_WBU_io_RegFileAccess_wd [2] ) );
BUF_X1 \WBU/_531_ ( .A(\_EXU_io_out_bits_memOut [3] ), .Z(\WBU/_126_ ) );
BUF_X1 \WBU/_532_ ( .A(\_EXU_io_out_bits_aluOut [3] ), .Z(\WBU/_058_ ) );
BUF_X1 \WBU/_533_ ( .A(\WBU/_025_ ), .Z(\_WBU_io_RegFileAccess_wd [3] ) );
BUF_X1 \WBU/_534_ ( .A(\_EXU_io_out_bits_memOut [4] ), .Z(\WBU/_127_ ) );
BUF_X1 \WBU/_535_ ( .A(\_EXU_io_out_bits_aluOut [4] ), .Z(\WBU/_059_ ) );
BUF_X1 \WBU/_536_ ( .A(\WBU/_026_ ), .Z(\_WBU_io_RegFileAccess_wd [4] ) );
BUF_X1 \WBU/_537_ ( .A(\_EXU_io_out_bits_memOut [5] ), .Z(\WBU/_128_ ) );
BUF_X1 \WBU/_538_ ( .A(\_EXU_io_out_bits_aluOut [5] ), .Z(\WBU/_060_ ) );
BUF_X1 \WBU/_539_ ( .A(\WBU/_027_ ), .Z(\_WBU_io_RegFileAccess_wd [5] ) );
BUF_X1 \WBU/_540_ ( .A(\_EXU_io_out_bits_memOut [6] ), .Z(\WBU/_129_ ) );
BUF_X1 \WBU/_541_ ( .A(\_EXU_io_out_bits_aluOut [6] ), .Z(\WBU/_061_ ) );
BUF_X1 \WBU/_542_ ( .A(\WBU/_028_ ), .Z(\_WBU_io_RegFileAccess_wd [6] ) );
BUF_X1 \WBU/_543_ ( .A(\_EXU_io_out_bits_memOut [7] ), .Z(\WBU/_130_ ) );
BUF_X1 \WBU/_544_ ( .A(\_EXU_io_out_bits_aluOut [7] ), .Z(\WBU/_062_ ) );
BUF_X1 \WBU/_545_ ( .A(\WBU/_029_ ), .Z(\_WBU_io_RegFileAccess_wd [7] ) );
BUF_X1 \WBU/_546_ ( .A(\_EXU_io_out_bits_memOut [8] ), .Z(\WBU/_131_ ) );
BUF_X1 \WBU/_547_ ( .A(\_EXU_io_out_bits_aluOut [8] ), .Z(\WBU/_063_ ) );
BUF_X1 \WBU/_548_ ( .A(\WBU/_030_ ), .Z(\_WBU_io_RegFileAccess_wd [8] ) );
BUF_X1 \WBU/_549_ ( .A(\_EXU_io_out_bits_memOut [9] ), .Z(\WBU/_132_ ) );
BUF_X1 \WBU/_550_ ( .A(\_EXU_io_out_bits_aluOut [9] ), .Z(\WBU/_064_ ) );
BUF_X1 \WBU/_551_ ( .A(\WBU/_031_ ), .Z(\_WBU_io_RegFileAccess_wd [9] ) );
BUF_X1 \WBU/_552_ ( .A(\_EXU_io_out_bits_memOut [10] ), .Z(\WBU/_102_ ) );
BUF_X1 \WBU/_553_ ( .A(\_EXU_io_out_bits_aluOut [10] ), .Z(\WBU/_034_ ) );
BUF_X1 \WBU/_554_ ( .A(\WBU/_001_ ), .Z(\_WBU_io_RegFileAccess_wd [10] ) );
BUF_X1 \WBU/_555_ ( .A(\_EXU_io_out_bits_memOut [11] ), .Z(\WBU/_103_ ) );
BUF_X1 \WBU/_556_ ( .A(\_EXU_io_out_bits_aluOut [11] ), .Z(\WBU/_035_ ) );
BUF_X1 \WBU/_557_ ( .A(\WBU/_002_ ), .Z(\_WBU_io_RegFileAccess_wd [11] ) );
BUF_X1 \WBU/_558_ ( .A(\_EXU_io_out_bits_memOut [12] ), .Z(\WBU/_104_ ) );
BUF_X1 \WBU/_559_ ( .A(\_EXU_io_out_bits_aluOut [12] ), .Z(\WBU/_036_ ) );
BUF_X1 \WBU/_560_ ( .A(\WBU/_003_ ), .Z(\_WBU_io_RegFileAccess_wd [12] ) );
BUF_X1 \WBU/_561_ ( .A(\_EXU_io_out_bits_memOut [13] ), .Z(\WBU/_105_ ) );
BUF_X1 \WBU/_562_ ( .A(\_EXU_io_out_bits_aluOut [13] ), .Z(\WBU/_037_ ) );
BUF_X1 \WBU/_563_ ( .A(\WBU/_004_ ), .Z(\_WBU_io_RegFileAccess_wd [13] ) );
BUF_X1 \WBU/_564_ ( .A(\_EXU_io_out_bits_memOut [14] ), .Z(\WBU/_106_ ) );
BUF_X1 \WBU/_565_ ( .A(\_EXU_io_out_bits_aluOut [14] ), .Z(\WBU/_038_ ) );
BUF_X1 \WBU/_566_ ( .A(\WBU/_005_ ), .Z(\_WBU_io_RegFileAccess_wd [14] ) );
BUF_X1 \WBU/_567_ ( .A(\_EXU_io_out_bits_memOut [15] ), .Z(\WBU/_107_ ) );
BUF_X1 \WBU/_568_ ( .A(\_EXU_io_out_bits_aluOut [15] ), .Z(\WBU/_039_ ) );
BUF_X1 \WBU/_569_ ( .A(\WBU/_006_ ), .Z(\_WBU_io_RegFileAccess_wd [15] ) );
BUF_X1 \WBU/_570_ ( .A(\_EXU_io_out_bits_memOut [16] ), .Z(\WBU/_108_ ) );
BUF_X1 \WBU/_571_ ( .A(\_EXU_io_out_bits_aluOut [16] ), .Z(\WBU/_040_ ) );
BUF_X1 \WBU/_572_ ( .A(\WBU/_007_ ), .Z(\_WBU_io_RegFileAccess_wd [16] ) );
BUF_X1 \WBU/_573_ ( .A(\_EXU_io_out_bits_memOut [17] ), .Z(\WBU/_109_ ) );
BUF_X1 \WBU/_574_ ( .A(\_EXU_io_out_bits_aluOut [17] ), .Z(\WBU/_041_ ) );
BUF_X1 \WBU/_575_ ( .A(\WBU/_008_ ), .Z(\_WBU_io_RegFileAccess_wd [17] ) );
BUF_X1 \WBU/_576_ ( .A(\_EXU_io_out_bits_memOut [18] ), .Z(\WBU/_110_ ) );
BUF_X1 \WBU/_577_ ( .A(\_EXU_io_out_bits_aluOut [18] ), .Z(\WBU/_042_ ) );
BUF_X1 \WBU/_578_ ( .A(\WBU/_009_ ), .Z(\_WBU_io_RegFileAccess_wd [18] ) );
BUF_X1 \WBU/_579_ ( .A(\_EXU_io_out_bits_memOut [19] ), .Z(\WBU/_111_ ) );
BUF_X1 \WBU/_580_ ( .A(\_EXU_io_out_bits_aluOut [19] ), .Z(\WBU/_043_ ) );
BUF_X1 \WBU/_581_ ( .A(\WBU/_010_ ), .Z(\_WBU_io_RegFileAccess_wd [19] ) );
BUF_X1 \WBU/_582_ ( .A(\_EXU_io_out_bits_memOut [20] ), .Z(\WBU/_113_ ) );
BUF_X1 \WBU/_583_ ( .A(\_EXU_io_out_bits_aluOut [20] ), .Z(\WBU/_045_ ) );
BUF_X1 \WBU/_584_ ( .A(\WBU/_012_ ), .Z(\_WBU_io_RegFileAccess_wd [20] ) );
BUF_X1 \WBU/_585_ ( .A(\_EXU_io_out_bits_memOut [21] ), .Z(\WBU/_114_ ) );
BUF_X1 \WBU/_586_ ( .A(\_EXU_io_out_bits_aluOut [21] ), .Z(\WBU/_046_ ) );
BUF_X1 \WBU/_587_ ( .A(\WBU/_013_ ), .Z(\_WBU_io_RegFileAccess_wd [21] ) );
BUF_X1 \WBU/_588_ ( .A(\_EXU_io_out_bits_memOut [22] ), .Z(\WBU/_115_ ) );
BUF_X1 \WBU/_589_ ( .A(\_EXU_io_out_bits_aluOut [22] ), .Z(\WBU/_047_ ) );
BUF_X1 \WBU/_590_ ( .A(\WBU/_014_ ), .Z(\_WBU_io_RegFileAccess_wd [22] ) );
BUF_X1 \WBU/_591_ ( .A(\_EXU_io_out_bits_memOut [23] ), .Z(\WBU/_116_ ) );
BUF_X1 \WBU/_592_ ( .A(\_EXU_io_out_bits_aluOut [23] ), .Z(\WBU/_048_ ) );
BUF_X1 \WBU/_593_ ( .A(\WBU/_015_ ), .Z(\_WBU_io_RegFileAccess_wd [23] ) );
BUF_X1 \WBU/_594_ ( .A(\_EXU_io_out_bits_memOut [24] ), .Z(\WBU/_117_ ) );
BUF_X1 \WBU/_595_ ( .A(\_EXU_io_out_bits_aluOut [24] ), .Z(\WBU/_049_ ) );
BUF_X1 \WBU/_596_ ( .A(\WBU/_016_ ), .Z(\_WBU_io_RegFileAccess_wd [24] ) );
BUF_X1 \WBU/_597_ ( .A(\_EXU_io_out_bits_memOut [25] ), .Z(\WBU/_118_ ) );
BUF_X1 \WBU/_598_ ( .A(\_EXU_io_out_bits_aluOut [25] ), .Z(\WBU/_050_ ) );
BUF_X1 \WBU/_599_ ( .A(\WBU/_017_ ), .Z(\_WBU_io_RegFileAccess_wd [25] ) );
BUF_X1 \WBU/_600_ ( .A(\_EXU_io_out_bits_memOut [26] ), .Z(\WBU/_119_ ) );
BUF_X1 \WBU/_601_ ( .A(\_EXU_io_out_bits_aluOut [26] ), .Z(\WBU/_051_ ) );
BUF_X1 \WBU/_602_ ( .A(\WBU/_018_ ), .Z(\_WBU_io_RegFileAccess_wd [26] ) );
BUF_X1 \WBU/_603_ ( .A(\_EXU_io_out_bits_memOut [27] ), .Z(\WBU/_120_ ) );
BUF_X1 \WBU/_604_ ( .A(\_EXU_io_out_bits_aluOut [27] ), .Z(\WBU/_052_ ) );
BUF_X1 \WBU/_605_ ( .A(\WBU/_019_ ), .Z(\_WBU_io_RegFileAccess_wd [27] ) );
BUF_X1 \WBU/_606_ ( .A(\_EXU_io_out_bits_memOut [28] ), .Z(\WBU/_121_ ) );
BUF_X1 \WBU/_607_ ( .A(\_EXU_io_out_bits_aluOut [28] ), .Z(\WBU/_053_ ) );
BUF_X1 \WBU/_608_ ( .A(\WBU/_020_ ), .Z(\_WBU_io_RegFileAccess_wd [28] ) );
BUF_X1 \WBU/_609_ ( .A(\_EXU_io_out_bits_memOut [29] ), .Z(\WBU/_122_ ) );
BUF_X1 \WBU/_610_ ( .A(\_EXU_io_out_bits_aluOut [29] ), .Z(\WBU/_054_ ) );
BUF_X1 \WBU/_611_ ( .A(\WBU/_021_ ), .Z(\_WBU_io_RegFileAccess_wd [29] ) );
BUF_X1 \WBU/_612_ ( .A(\_EXU_io_out_bits_memOut [30] ), .Z(\WBU/_124_ ) );
BUF_X1 \WBU/_613_ ( .A(\_EXU_io_out_bits_aluOut [30] ), .Z(\WBU/_056_ ) );
BUF_X1 \WBU/_614_ ( .A(\WBU/_023_ ), .Z(\_WBU_io_RegFileAccess_wd [30] ) );
BUF_X1 \WBU/_615_ ( .A(\_EXU_io_out_bits_memOut [31] ), .Z(\WBU/_125_ ) );
BUF_X1 \WBU/_616_ ( .A(\_EXU_io_out_bits_aluOut [31] ), .Z(\WBU/_057_ ) );
BUF_X1 \WBU/_617_ ( .A(\WBU/_024_ ), .Z(\_WBU_io_RegFileAccess_wd [31] ) );
BUF_X1 \WBU/_618_ ( .A(_EXU_io_out_valid ), .Z(\WBU/_165_ ) );
BUF_X1 \WBU/_619_ ( .A(_EXU_io_out_bits_control_regWe ), .Z(\WBU/_066_ ) );
BUF_X1 \WBU/_620_ ( .A(\WBU/_032_ ), .Z(_WBU_io_RegFileAccess_we ) );
BUF_X8 fanout_buf_1 ( .A(_00_ ), .Z(fanout_net_1 ) );
BUF_X8 fanout_buf_2 ( .A(_00_ ), .Z(fanout_net_2 ) );
BUF_X8 fanout_buf_3 ( .A(\AXI4Interconnect/_0004_ ), .Z(fanout_net_3 ) );
BUF_X8 fanout_buf_4 ( .A(\AXI4Interconnect/_0004_ ), .Z(fanout_net_4 ) );
BUF_X8 fanout_buf_5 ( .A(\AXI4Interconnect/_0869_ ), .Z(fanout_net_5 ) );
BUF_X8 fanout_buf_6 ( .A(\AXI4Interconnect/_0871_ ), .Z(fanout_net_6 ) );
BUF_X8 fanout_buf_7 ( .A(\CLINT/_0577_ ), .Z(fanout_net_7 ) );
BUF_X8 fanout_buf_8 ( .A(\EXU/_0067_ ), .Z(fanout_net_8 ) );
BUF_X8 fanout_buf_9 ( .A(\EXU/_0068_ ), .Z(fanout_net_9 ) );
BUF_X8 fanout_buf_10 ( .A(\EXU/_0381_ ), .Z(fanout_net_10 ) );
BUF_X8 fanout_buf_11 ( .A(\EXU/_0394_ ), .Z(fanout_net_11 ) );
BUF_X8 fanout_buf_12 ( .A(\EXU/ALU/_034_ ), .Z(fanout_net_12 ) );
BUF_X8 fanout_buf_13 ( .A(\EXU/ALU/_035_ ), .Z(fanout_net_13 ) );
BUF_X8 fanout_buf_14 ( .A(\EXU/ALU/_036_ ), .Z(fanout_net_14 ) );
BUF_X8 fanout_buf_15 ( .A(\EXU/ALU/_036_ ), .Z(fanout_net_15 ) );
BUF_X8 fanout_buf_16 ( .A(\EXU/ALU/adder/_000_ ), .Z(fanout_net_16 ) );
BUF_X8 fanout_buf_17 ( .A(\EXU/CSRControl/_0272_ ), .Z(fanout_net_17 ) );
BUF_X8 fanout_buf_18 ( .A(\EXU/CSRControl/_0273_ ), .Z(fanout_net_18 ) );
BUF_X8 fanout_buf_19 ( .A(\LSU/_0316_ ), .Z(fanout_net_19 ) );
BUF_X8 fanout_buf_20 ( .A(\WBU/_065_ ), .Z(fanout_net_20 ) );

endmodule
